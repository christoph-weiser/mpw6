* SPICE3 file created from main.ext - technology: sky130A


.subckt main dvdd en_ldo_dig avdd rstn vdd vss en_ldo_ana clksys en_clk_int clkext ibp_3_ ibp_2_
+ ibp_1_ ibp_0_ ibn_1_ ibn_0_ en_clkdiv clksel refsel vbg_ext avss dvss tbout bgtrim_15_ bgtrim_14_
+ bgtrim_13_ bgtrim_12_ bgtrim_11_ bgtrim_10_ bgtrim_9_ bgtrim_8_ bgtrim_7_ bgtrim_6_ bgtrim_5_ bgtrim_4_
+ bgtrim_3_ bgtrim_2_ bgtrim_1_ bgtrim_0_ tbctl_2_ tbctl_1_ tbctl_0_

Rconn1 avss vss 0.01
Rconn2 dvss vss 0.01

X0 a_29435_30536# a_30910_30664# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=9.28e+12p pd=8.256e+07u as=9.28e+12p ps=8.256e+07u w=1e+06u l=500000u
X2 a_16019_26544# a_7257_35054# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=1.032e+07u as=4.64e+12p ps=4.128e+07u w=1e+06u l=4e+06u
X3 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.42759e+14p pd=2.04143e+09u as=0p ps=0u w=870000u l=1.05e+06u
X4 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.66245e+14p pd=1.47076e+09u as=0p ps=0u w=2e+06u l=4e+06u
X5 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X6 a_21533_59718# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=6.38e+12p pd=5.676e+07u as=0p ps=0u w=1e+06u l=1e+06u
X7 a_27549_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=2.064e+07u as=4.582e+13p ps=3.3862e+08u w=1e+06u l=1e+06u
X8 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X9 vss ibp_2_ ibp_2_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.61e+12p ps=2.322e+07u w=1e+06u l=1e+06u
X10 a_8302_16888# a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.61e+12p pd=2.322e+07u as=0p ps=0u w=1e+06u l=500000u
X11 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X12 a_39286_5164# a_38770_5164# a_39191_5164# vss sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X13 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X14 a_17509_48421# a_17233_48421# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X15 vss ibpbas a_16196_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=6.32e+06u w=500000u l=4e+06u
X16 vdd a_14147_17413# a_23557_19518# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X17 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X18 vdd a_10803_51693# a_8735_54512# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X19 a_9785_4482# ibp_1_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=4.64e+12p pd=4.128e+07u as=0p ps=0u w=1e+06u l=1e+06u
X20 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.624e+13p ps=1.352e+08u w=1e+06u l=1e+06u
X21 a_21272_47107# ibp_0_ ibp_0_ vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.406e+07u as=1.16e+12p ps=9.16e+06u w=2e+06u l=4e+06u
X22 a_9727_51399# a_9697_51123# a_9473_51399# vdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X23 a_46660_5972# a_46036_5606# a_46552_5606# dvdd sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X24 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X25 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X26 a_47409_7016# a_46031_4206# a_46897_6668# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.344e+11p pd=1.7e+06u as=2.624e+11p ps=2.1e+06u w=640000u l=150000u
X27 a_28184_49195# a_28184_49195# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=4.06e+12p pd=3.612e+07u as=6.38e+12p ps=5.676e+07u w=1e+06u l=4e+06u
X28 dvdd a_46031_5294# a_46036_5068# dvdd sky130_fd_pr__pfet_01v8_hvt ad=5.7007e+13p pd=4.5023e+08u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X29 a_29435_33716# bgtrim_8_ a_29277_29476# vss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=9.28e+12p ps=7.328e+07u w=2e+06u l=500000u
X30 vdd en_ldo_dig a_40013_15426# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.548e+07u w=1e+06u l=400000u
X31 dvdd a_46031_4206# a_46036_3980# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X32 ibp_2_ ibp_2_ ibp_2_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X33 vss a_9183_51693# a_10895_50605# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X34 a_21333_59018# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X35 dvdd a_46770_5848# a_46660_5972# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_8735_54512# a_10803_51693# vss vss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X37 a_29435_36896# a_30910_37024# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X38 vbg a_7028_39565# vbg_ext vdd sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X39 a_9039_52781# a_8871_52781# vss vss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X40 ibp_2_ ibp_2_ vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X41 a_16019_27456# ibnbas a_15161_31718# vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=1.832e+07u as=9.28e+12p ps=7.328e+07u w=2e+06u l=4e+06u
X42 a_6633_29468# a_6949_30834# a_7149_30931# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.827e+13p pd=1.3818e+08u as=4.64e+12p ps=3.432e+07u w=4e+06u l=1e+06u
X43 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X44 a_14147_17413# a_14147_17185# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=6.32e+06u as=0p ps=0u w=500000u l=1e+07u
X45 a_7149_30931# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=4.64e+12p pd=4.128e+07u as=0p ps=0u w=1e+06u l=1e+06u
X46 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X47 vbg a_8742_39565# vbg_int vss sky130_fd_pr__nfet_01v8 ad=8.7e+11p pd=7.74e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X48 a_27033_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=4.64e+12p pd=4.128e+07u as=0p ps=0u w=1e+06u l=1e+06u
X49 a_36712_33396# a_36326_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X50 vss a_27549_7238# a_27549_7238# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.548e+07u w=1e+06u l=1e+06u
X51 a_7257_35054# a_7257_35054# a_7257_35054# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.58e+07u as=0p ps=0u w=1e+06u l=4e+06u
X52 vss a_6880_26619# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X53 a_14147_17413# a_14605_15614# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X54 vdd a_8735_54512# a_10773_52781# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X55 a_10533_55475# a_8735_54512# vss vss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X56 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X57 a_9340_13770# vss vss sky130_fd_pr__res_xhigh_po w=350000u l=7e+06u
X58 a_9033_7909# en_ldo_ana vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.548e+07u as=0p ps=0u w=1e+06u l=400000u
X59 a_16019_26544# ibnbas a_15161_30727# vdd sky130_fd_pr__pfet_01v8_lvt ad=6.96e+12p pd=5.496e+07u as=9.28e+12p ps=7.328e+07u w=2e+06u l=4e+06u
X60 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.624e+13p pd=1.352e+08u as=0p ps=0u w=1e+06u l=1e+06u
X61 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X62 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X63 vdd a_16019_26544# a_15161_30727# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X64 a_39504_5406# a_39286_5164# vss vss sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X65 vss a_10117_54413# a_10283_54413# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X66 a_29277_29476# bgtrim_13_ a_30910_35964# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X67 a_46770_4760# a_46552_4518# vss vss sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X68 a_9785_4482# ibp_1_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X69 vdd a_21333_59018# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X70 vss ibp_1_ ibp_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.61e+12p ps=2.322e+07u w=1e+06u l=1e+06u
X71 avdd a_9033_7909# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X72 a_29267_5405# a_27549_7238# vss vss sky130_fd_pr__nfet_01v8 ad=3.19e+12p pd=2.838e+07u as=0p ps=0u w=1e+06u l=1e+06u
X73 vss a_27549_7238# a_27549_7238# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X74 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X75 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X76 a_9371_53985# a_8861_54387# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X77 vss a_21272_47107# a_21088_54984# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=1.032e+07u w=1e+06u l=1e+06u
X78 vdd a_10803_51693# a_8735_54512# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X79 vdd a_16019_26544# a_15161_30727# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X80 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X81 vdd a_10287_50605# a_11129_51149# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X82 a_21030_55081# a_21088_54984# a_21088_54984# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.29e+07u as=5.8e+11p ps=5.16e+06u w=1e+06u l=4e+06u
X83 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X84 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X85 a_16534_48421# a_16071_51406# dvdd vss sky130_fd_pr__nfet_01v8 ad=2.32e+12p pd=2.064e+07u as=1.04237e+13p ps=1.2588e+08u w=1e+06u l=500000u
X86 a_21230_16137# a_21230_16137# a_22146_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=1.16e+12p ps=1.032e+07u w=1e+06u l=2e+06u
X87 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X88 vdd a_21030_55081# a_21030_55081# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X89 tbout a_28184_48339# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=3.48e+12p pd=2.574e+07u as=0p ps=0u w=4e+06u l=4e+06u
X90 a_28184_48339# a_28184_48339# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=4.06e+12p pd=3.612e+07u as=0p ps=0u w=1e+06u l=4e+06u
X91 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X92 a_9033_6762# en_ldo_ana vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X93 a_43124_15781# a_37846_16790# a_40013_15754# vss sky130_fd_pr__nfet_01v8_lvt ad=4.64e+12p pd=4.128e+07u as=2.03e+12p ps=1.806e+07u w=1e+06u l=1e+06u
X94 a_22146_16137# a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X95 a_11221_50213# a_11129_51149# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X96 avdd a_9033_7909# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X97 a_46247_6846# clksel vss vss sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X98 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X99 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X100 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X101 vdd a_11221_50061# a_11398_50061# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X102 a_16534_48421# a_16071_57376# avdd vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.75807e+13p ps=2.06e+08u w=1e+06u l=500000u
X103 ibp_2_ ibp_2_ ibp_2_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X104 a_16071_54391# a_15795_54391# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X105 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X106 vdd a_21333_59018# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X107 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X108 a_47279_3974# a_46202_3980# a_47117_4352# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X109 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X110 a_21257_48618# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.044e+13p pd=8.476e+07u as=0p ps=0u w=1e+06u l=1e+06u
X111 a_21533_59718# a_16534_48421# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.832e+07u as=0p ps=0u w=2e+06u l=1e+06u
X112 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X113 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X114 vdd a_9091_54413# a_9473_54965# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X115 a_21015_51763# a_16534_48421# a_21531_53226# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.856e+13p pd=1.4076e+08u as=4.64e+12p ps=3.432e+07u w=4e+06u l=1e+06u
X116 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X117 vb_6_ a_32117_14563# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X118 a_7973_17910# a_7973_17910# a_7909_15880# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+11p pd=1.58e+06u as=1.45e+11p ps=1.58e+06u w=500000u l=1e+06u
X119 a_29435_33716# a_30910_32784# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X120 a_17146_5558# a_16724_7690# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X121 vss a_9697_51123# a_9521_52211# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X122 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X123 vdd a_14147_17413# a_14605_15614# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=1.264e+07u w=500000u l=2e+06u
R0 vss vss sky130_fd_pr__res_generic_m4 w=9.6e+06u l=4e+06u
X124 a_21333_59018# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X125 a_48035_5606# a_47856_5606# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X126 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X127 a_21531_51763# ibp_0_ a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.12e+12p ps=6.412e+07u w=2e+06u l=4e+06u
X128 vdd a_21333_59018# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X129 a_21531_51763# ibp_0_ a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X130 a_16019_27456# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X131 a_7057_34366# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.432e+07u as=0p ps=0u w=1e+06u l=1e+06u
X132 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X133 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X134 a_46340_4145# a_46031_4670# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X135 a_7257_35054# a_7257_35054# a_7257_35054# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X136 a_21257_48618# a_16534_48421# a_21533_59718# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X137 vdd a_8871_56045# a_8933_54387# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X138 a_8819_54413# a_8735_54512# a_8737_54413# vss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X139 w_42506_30499# w_42506_30499# vdd vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=1e+06u
X140 a_16534_48421# a_17509_51406# vb_4_ vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X141 a_17509_54391# a_17233_54391# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X142 a_8302_16888# a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X143 a_21793_20190# a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=0p ps=0u w=500000u l=2e+06u
X144 vdd a_21030_55081# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X145 vss ibp_2_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X146 vss a_10197_55475# a_10227_55501# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X147 a_8302_16888# a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=0p ps=0u w=1e+06u l=1e+06u
X148 vdd a_14147_17413# a_14605_15614# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X149 vss a_6880_26619# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X150 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X151 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X152 a_9567_53869# a_8735_54512# vss vss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X153 a_33084_6373# a_33004_6347# a_29267_5405# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X154 vdd a_14147_17413# a_14605_15614# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X155 a_33004_6347# a_35079_6373# a_29267_5405# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X156 a_16534_48421# a_17509_57376# vdd vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.61908e+14p ps=3.08131e+09u w=1e+06u l=500000u
X157 avdd ibn_0_ a_27549_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X158 a_7080_26645# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X159 a_11926_4549# a_12242_4494# a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=2.03e+12p pd=1.806e+07u as=0p ps=0u w=1e+06u l=1e+06u
X160 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X161 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X162 vdd a_9105_50837# a_9105_50605# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X163 vss a_9013_51925# a_9013_51693# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X164 a_9091_54413# a_8737_54413# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X165 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X166 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X167 a_10073_52389# a_10346_52217# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X168 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X169 a_47292_4278# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X170 vdd a_7057_34366# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X171 a_28184_48339# ibp_0_ a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=8.12e+12p pd=6.412e+07u as=0p ps=0u w=2e+06u l=4e+06u
X172 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X173 ibn_1_ a_21230_16137# ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=0p ps=0u w=1e+06u l=2e+06u
X174 ibn_1_ a_21230_16137# a_23062_17193# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X175 dvdd a_47292_4278# a_47856_3974# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X176 a_7080_26645# a_6949_29442# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.432e+07u as=0p ps=0u w=4e+06u l=1e+06u
X177 vss a_21230_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X178 ibpbas a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=1e+06u
X179 a_23062_17193# a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X180 a_15161_30727# ibnbas a_16019_26544# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X181 a_9936_52053# a_9039_52781# a_9855_52053# vss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X182 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X183 vb_0_ a_32117_20471# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X184 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X185 a_16196_13967# ibpbas a_15338_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=1.264e+07u w=500000u l=4e+06u
X186 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X187 vss a_10895_50605# a_11063_50605# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X188 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X189 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X190 ibnbas a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=500000u
X191 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X192 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X193 a_10383_52897# a_9697_51123# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X194 a_14147_17413# a_14605_15614# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X195 a_10018_50965# a_9831_50605# a_9931_50721# vss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X196 a_9785_4482# a_12242_4494# a_11926_4549# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X197 a_15161_31718# ibnbas a_16019_27456# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X198 vss a_10117_54413# a_10283_54413# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X199 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X200 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X201 vss a_47292_5580# a_47856_5606# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X202 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X203 a_10073_52389# a_10346_52217# a_10304_52243# vss sky130_fd_pr__nfet_01v8 ad=1.07825e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X204 vss a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X205 a_28184_48339# a_28184_49195# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X206 avdd ibn_0_ a_27033_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X207 vss a_21230_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X208 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X209 a_8735_54512# a_10803_51693# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X210 a_21531_51763# ibp_0_ a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X211 a_47117_4518# a_46036_4518# a_46770_4760# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X212 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X213 a_10533_56019# a_9697_51123# a_10593_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=7.9e+11p ps=7.58e+06u w=1e+06u l=150000u
X214 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X215 a_9785_4482# a_12242_4494# a_11926_4549# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X216 vss a_6880_26619# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X217 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X218 vss a_10143_50061# a_17233_48421# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X219 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X220 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X221 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X222 a_46552_5440# a_46202_5068# a_46457_5428# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X223 vss a_47292_4278# a_47226_4352# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X224 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X225 a_21531_53226# ibp_0_ a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X226 a_11398_50061# a_11221_50061# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X227 a_21333_59018# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X228 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X229 a_27549_7238# a_27549_7238# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X230 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X231 vdd a_7057_34366# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X232 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X233 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X234 a_37846_16790# a_37846_18922# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X235 a_39548_5164# a_39504_5406# a_39382_5164# vss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X236 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X237 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X238 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X239 a_21533_59718# a_16534_48421# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X240 a_16019_26544# a_7257_35054# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X241 a_27549_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X242 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X243 a_34723_6373# a_34367_6373# a_27033_7238# avdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X244 vdd a_7057_34366# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X245 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X246 a_21015_51763# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X247 a_8302_16888# a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X248 avdd ibn_0_ a_27549_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X249 vdd a_9506_17973# a_8302_16888# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X250 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X251 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X252 a_40013_15754# a_40013_15754# a_40013_15754# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X253 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X254 a_28184_48339# ibp_0_ a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X255 a_10287_50605# a_9931_50721# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X256 vss a_16302_7690# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X257 a_29435_31596# bgtrim_4_ a_29277_29476# vss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X258 a_47471_4340# rstn vss vss sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X259 ibnbas ibnbas ibnbas vdd sky130_fd_pr__pfet_01v8_lvt ad=6.96e+12p pd=5.496e+07u as=0p ps=0u w=2e+06u l=4e+06u
X260 ibpbas ibpbas vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=1.264e+07u as=0p ps=0u w=500000u l=4e+06u
X261 vdd a_10435_54957# a_9697_51123# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X262 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X263 ibp_1_ a_14147_17413# a_21793_19294# vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X264 vdd a_7057_34366# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X265 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X266 vss a_9977_51123# a_9521_52211# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X267 a_16534_48421# a_15795_57376# avdd vdd sky130_fd_pr__pfet_01v8 ad=2.32e+12p pd=2.064e+07u as=0p ps=0u w=1e+06u l=500000u
X268 a_33084_7058# vss sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=4e+06u
X269 a_21531_53226# a_16534_48421# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X270 a_9033_6762# en_ldo_ana vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X271 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X272 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X273 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X274 a_46897_6668# a_47267_6832# a_47124_7016# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.576e+11p ps=2.71e+06u w=640000u l=150000u
X275 a_6633_29468# a_6949_30834# a_7149_30931# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X276 dvdd a_40013_15426# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X277 vss rstn a_46814_4340# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X278 ibnbas ibnbas ibnbas vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X279 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X280 vdd a_9506_17973# ibpbas vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X281 a_16196_13967# ibpbas vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X282 vb_2_ a_32117_18783# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X283 a_21531_53226# a_16534_48421# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X284 a_9521_52211# a_9697_51123# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X285 vss a_47292_5366# a_47856_5062# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X286 a_9033_7909# a_11926_4549# a_9033_7909# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X287 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X288 a_46770_4760# a_46552_4518# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X289 a_28184_48339# a_28184_49195# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X290 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X291 a_14147_17185# a_14147_17185# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=6.32e+06u as=0p ps=0u w=500000u l=1e+07u
X292 a_28184_48339# ibp_0_ a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X293 vss a_10803_51693# a_8735_54512# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X294 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X295 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X296 a_21533_59718# a_16534_48421# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X297 vdd a_9697_51123# a_10073_52389# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X298 a_37098_33396# a_35940_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X299 dvdd a_47117_4518# a_47292_4492# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X300 a_9785_4482# ibp_1_ vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X301 vss a_46031_4206# a_46036_3980# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X302 avdd ibn_0_ a_27549_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X303 a_28184_48339# a_28184_49195# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X304 dvdd clksel a_46581_7016# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.344e+11p ps=1.7e+06u w=640000u l=150000u
X305 a_7149_30931# a_7257_35054# a_16019_27456# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+12p ps=1.29e+07u w=1e+06u l=4e+06u
X306 vdd a_11398_50061# a_15795_48421# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X307 vss a_10895_50605# a_11063_50605# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X308 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X309 vss a_9065_53299# a_8861_54387# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X310 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X311 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X312 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X313 a_21531_53226# ibp_0_ a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X314 vss tbctl_2_ a_8737_50061# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X315 avdd ibn_0_ a_27549_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X316 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X317 a_9506_17973# a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=0p ps=0u w=1e+06u l=1e+06u
X318 a_21333_59018# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X319 vss a_47292_4492# a_47226_4518# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.338e+11p ps=1.5e+06u w=420000u l=150000u
X320 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X321 vss a_47886_16107# ibp_2_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=400000u
X322 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X323 a_16534_48421# a_17233_57376# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X324 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X325 a_10865_53869# a_8861_54387# a_10593_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u
X326 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X327 a_16019_27456# a_7257_35054# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X328 a_7080_26645# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X329 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X330 vdd a_40013_15754# a_40013_15754# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.45e+12p ps=1.29e+07u w=1e+06u l=1e+06u
X331 a_21257_48618# a_16534_48421# a_21533_59718# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X332 vss vss a_29277_29476# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=3.6992e+12p
X333 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X334 a_21531_51763# tbout a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=4.64e+12p pd=3.432e+07u as=0p ps=0u w=4e+06u l=1e+06u
X335 a_29435_34776# bgtrim_10_ a_29277_29476# vss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X336 a_8302_16888# a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X337 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X338 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X339 a_6633_29468# a_6633_29468# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X340 a_10533_56019# a_8861_54387# vss vss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X341 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X342 a_39851_5164# a_38770_5164# a_39504_5406# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X343 a_46340_5819# a_47267_6832# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X344 a_47279_5972# a_46202_5606# a_47117_5606# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X345 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X346 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X347 dvdd a_46927_6694# a_47756_6694# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.8e+11p ps=2.56e+06u w=1e+06u l=150000u
X348 a_8302_16888# a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X349 vss a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X350 a_39504_5406# a_39286_5164# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X351 a_47267_6832# a_47292_5580# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X352 a_11926_4549# a_11926_4549# a_11926_4549# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.29e+07u as=0p ps=0u w=1e+06u l=1e+06u
X353 a_46340_4731# a_46031_5294# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X354 a_47471_4518# rstn vss vss sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X355 a_8302_16888# a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X356 vss a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X357 a_46660_3974# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X358 avdd ibn_0_ a_27033_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X359 a_9785_4482# ibp_1_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X360 a_27033_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X361 vss a_11398_53325# a_17233_54391# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X362 a_6880_26619# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.74e+12p pd=1.548e+07u as=0p ps=0u w=1e+06u l=1e+06u
X363 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X364 a_39382_5164# a_38936_5164# a_39286_5164# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X365 vdd a_11926_4549# a_9033_7909# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X366 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X367 a_28184_48339# a_28184_49195# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X368 vss a_46069_6668# a_46031_4206# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X369 a_11926_4549# a_11926_4549# a_11926_4549# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X370 a_48035_5062# a_47856_5062# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X371 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X372 vss a_28184_48339# tbout vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.48e+12p ps=2.574e+07u w=4e+06u l=4e+06u
X373 a_29277_29476# bgtrim_15_ a_30910_37024# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X374 a_10143_50061# a_9975_50061# vss vss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X375 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X376 a_10593_53869# a_8861_54387# a_10865_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X377 vss a_21230_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X378 vss rstn a_46814_4518# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X379 a_21272_47107# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X380 a_46457_5428# a_46340_5233# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X381 vss a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X382 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X383 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X384 a_28184_49195# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X385 a_23557_19518# a_14147_17413# a_21230_16137# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X386 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X387 a_46581_7016# a_40581_5164# a_46069_6668# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.624e+11p ps=2.1e+06u w=640000u l=150000u
X388 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X389 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X390 a_35079_6373# a_34723_6373# a_27033_7238# avdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X391 vdd a_40013_15754# a_40013_15426# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X392 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X393 vss ibp_1_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X394 a_29277_29476# bgtrim_1_ a_30910_29604# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X395 a_21230_16137# a_21230_16137# a_21230_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X396 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X397 dvdd a_40013_15426# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X398 vss vss a_6949_30834# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=4.624e+11p
X399 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X400 vdd a_14147_17185# a_14147_17185# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X401 ibp_0_ a_14147_17413# a_21793_19742# vdd sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=6.32e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X402 vdd a_16019_26544# a_15161_30727# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X403 a_27549_7238# a_27549_7238# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X404 a_28184_48339# a_28184_49195# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X405 vss a_46031_4670# a_46036_4518# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X406 vdd a_6416_39560# a_7028_39565# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X407 a_28184_48339# ibp_0_ a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X408 a_28184_48339# ibp_0_ a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X409 a_7080_26645# a_7257_35054# a_16019_26544# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X410 a_15161_31718# ibnbas a_16019_27456# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X411 a_9705_51925# a_8933_54387# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X412 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X413 a_47292_5580# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X414 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X415 a_43124_15781# vb_3_ a_40013_15426# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.03e+12p ps=1.806e+07u w=1e+06u l=1e+06u
X416 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X417 vss a_22146_16137# a_22146_15433# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X418 a_21257_48618# a_21257_48618# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X419 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X420 a_47396_6694# a_47267_6832# a_46897_6668# vss sky130_fd_pr__nfet_01v8 ad=1.155e+11p pd=1.39e+06u as=3.465e+11p ps=2.49e+06u w=420000u l=150000u
X421 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X422 a_22146_15433# a_21230_16137# ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X423 a_27033_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X424 a_9033_7909# vb_2_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=2.03e+12p pd=1.806e+07u as=0p ps=0u w=1e+06u l=1e+06u
R1 vss vss sky130_fd_pr__res_generic_m4 w=9.6e+06u l=4e+06u
X425 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X426 vdd a_16019_26544# a_15161_30727# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X427 a_8871_56045# tbctl_0_ vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X428 a_28184_48339# a_28184_48339# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X429 a_10593_53869# a_9697_51123# a_10533_56019# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X430 a_27549_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X431 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X432 a_15161_30727# ibnbas a_16019_26544# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X433 a_46278_6694# a_46247_6846# vss vss sky130_fd_pr__nfet_01v8 ad=1.365e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X434 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X435 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X436 vdd a_10227_55501# a_15795_57376# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X437 a_47292_5580# a_47117_5606# a_47471_5606# vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X438 a_33655_6373# vss sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=4e+06u
X439 a_16071_48421# a_15795_48421# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X440 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X441 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X442 ibp_0_ a_14147_17413# a_21793_19966# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X443 a_21533_59718# a_28184_49195# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X444 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X445 a_21015_51763# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X446 vss a_9105_50837# a_9105_50605# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X447 a_34723_6373# a_34367_6373# a_29267_5405# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X448 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X449 a_40205_5164# rstn vss vss sky130_fd_pr__nfet_01v8 ad=1.281e+11p pd=1.45e+06u as=0p ps=0u w=420000u l=150000u
X450 a_6633_29468# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X451 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X452 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X453 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X454 a_38936_5164# a_38770_5164# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X455 vss a_8861_54387# a_10533_55475# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X456 a_47075_6846# en_clkdiv dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.728e+11p pd=1.82e+06u as=0p ps=0u w=640000u l=150000u
X457 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X458 vss a_9039_52781# a_9065_53299# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X459 a_8861_54387# a_9065_53299# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X460 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X461 a_7149_30931# a_6949_30834# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X462 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X463 a_11063_50605# a_10895_50605# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X464 a_9785_4482# vb_2_ a_9033_7909# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X465 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X466 a_46660_4884# a_46036_4518# a_46552_4518# dvdd sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=1.449e+11p ps=1.53e+06u w=420000u l=150000u
X467 a_40572_33396# a_40958_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X468 a_16019_27456# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X469 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X470 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X471 vss a_21272_47107# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X472 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X473 vdd a_9506_17973# a_8302_16888# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X474 ibn_0_ ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=5.16e+06u as=0p ps=0u w=1e+06u l=1e+06u
X475 vss a_8735_54512# a_10533_55475# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X476 a_39851_5164# a_38936_5164# a_39504_5406# vss sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X477 a_15161_31718# a_16019_26544# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X478 vdd a_9065_53299# a_8861_54387# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X479 vdd a_16019_27456# a_39053_30692# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=1e+06u
X480 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X481 a_29435_33716# a_30910_33844# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X482 a_28184_49195# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X483 vdd tbctl_2_ a_8737_50061# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X484 a_21531_51763# ibp_0_ a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X485 a_7257_35054# a_7257_35054# a_6880_26619# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X486 a_28184_49195# a_28184_49195# a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X487 dvdd a_46770_4760# a_46660_4884# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X488 ibn_1_ a_21230_16137# ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X489 a_47117_4352# a_46202_3980# a_46770_3948# vss sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X490 vb_4_ a_32117_16251# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X491 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X492 a_38690_16790# a_39956_18922# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X493 vss vss vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X494 a_15161_31718# a_16019_26544# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X495 a_11063_50605# a_10895_50605# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X496 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X497 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X498 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X499 a_7909_13748# a_7909_15880# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X500 vss a_28184_48339# tbout vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X501 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X502 a_28184_48339# ibp_0_ a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X503 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X504 a_37098_33396# a_37484_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X505 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X506 a_10304_52243# a_9697_51123# a_10223_52243# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.071e+11p ps=1.35e+06u w=420000u l=150000u
X507 a_16019_27456# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X508 vdd a_14147_17413# a_14605_15614# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X509 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X510 vss ibpbas ibpbas vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X511 a_21533_59718# a_16534_48421# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X512 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X513 a_21015_51763# a_16534_48421# a_21531_53226# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X514 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X515 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X516 a_46552_4518# a_46036_4518# a_46457_4518# vss sky130_fd_pr__nfet_01v8 ad=1.188e+11p pd=1.38e+06u as=1.32e+11p ps=1.49e+06u w=360000u l=150000u
X517 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X518 a_47292_5366# a_47117_5440# a_47471_5428# vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=1.281e+11p ps=1.45e+06u w=420000u l=150000u
X519 a_48035_3974# a_47856_3974# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X520 a_21333_59018# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X521 a_40013_15426# vb_3_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X522 a_21257_48618# tbout a_21333_59018# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.32e+12p ps=1.832e+07u w=2e+06u l=1e+06u
X523 vss a_27549_7238# a_29267_5405# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X524 a_46202_5068# a_46036_5068# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X525 a_7304_39565# a_7028_39565# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X526 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X527 a_46202_3980# a_46036_3980# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X528 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X529 a_12242_4494# a_17990_7690# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X530 a_9727_51399# a_9977_51123# a_9521_52211# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X531 vss a_6880_26619# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X532 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X533 a_9215_52237# a_9185_52211# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X534 a_9506_17973# a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X535 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X536 a_34011_6373# a_33655_6373# a_27033_7238# avdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X537 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X538 vdd a_9039_52781# a_9065_53299# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X539 a_8121_17110# a_8121_17110# a_7973_17910# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+11p pd=1.58e+06u as=0p ps=0u w=500000u l=1e+06u
X540 vdd a_21030_55081# a_21030_55081# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X541 a_7080_26645# a_7257_35054# a_16019_26544# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X542 a_6880_26619# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X543 clksys a_47756_6694# vss vss sky130_fd_pr__nfet_01v8 ad=4.704e+11p pd=5.6e+06u as=0p ps=0u w=420000u l=150000u
X544 vdd a_14147_17413# a_23557_20190# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X545 a_9650_54957# a_9473_54965# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X546 vss a_9975_50061# a_10143_50061# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X547 vss a_9697_51123# a_9567_53869# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X548 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X549 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X550 a_14605_15614# a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X551 vdd a_8871_52781# a_9039_52781# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X552 a_47117_5606# a_46202_5606# a_46770_5848# vss sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=1.998e+11p ps=1.97e+06u w=360000u l=150000u
X553 a_21333_59018# tbout a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X554 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X555 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X556 a_7257_35054# a_7257_35054# a_6880_26619# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X557 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X558 a_21531_51763# ibp_0_ a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X559 a_48035_4518# a_47856_4518# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X560 vss refsel a_8466_39565# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X561 a_16071_54391# a_15795_54391# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X562 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X563 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X564 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X565 a_40013_15426# vb_3_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X566 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X567 a_35079_6373# a_34723_6373# a_29267_5405# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X568 a_46031_5758# a_47292_5366# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X569 dvdd a_40013_15426# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X570 a_8933_54387# a_8871_56045# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X571 a_8861_54387# a_9065_53299# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X572 a_11063_50605# a_10895_50605# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X573 a_21272_47107# ibp_0_ ibp_0_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X574 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X575 a_9033_7909# a_11926_4549# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X576 a_16019_26544# ibnbas a_15161_30727# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X577 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X578 a_15338_13967# ibpbas a_16196_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X579 a_9473_51399# a_8861_54387# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X580 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X581 a_28184_49195# a_28184_49195# a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X582 a_9215_52237# a_9185_52211# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X583 a_6633_29468# a_6949_29442# a_7080_26645# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X584 vdd a_21030_55081# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X585 a_40581_5164# a_40026_5138# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X586 a_48035_5606# a_47856_5606# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X587 a_8742_39565# a_8466_39565# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X588 a_46660_5972# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X589 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X590 a_8735_54512# a_10803_51693# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X591 a_28184_48339# a_28184_49195# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X592 a_39394_5530# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X593 a_21531_51763# tbout a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X594 a_17509_48421# a_17233_48421# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X595 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X596 dvdd a_47292_4278# a_47279_3974# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X597 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X598 a_16019_27456# ibnbas a_15161_31718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X599 vss a_47756_6694# clksys vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X600 vss ibpbas ibpbas vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X601 a_21333_59018# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X602 a_6949_29442# a_30910_37024# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X603 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X604 a_47124_7016# a_47075_6846# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X605 a_21257_48618# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X606 a_46814_5606# a_46770_5848# a_46648_5606# vss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X607 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X608 a_21533_59718# a_28184_49195# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X609 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X610 a_9065_53299# a_9039_52781# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X611 a_10533_55475# a_8861_54387# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X612 vdd tbctl_0_ a_8871_56045# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X613 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X614 vdd a_8871_52781# a_9039_52781# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X615 a_46897_6668# a_46031_4206# a_47106_6694# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=150000u
X616 a_10773_52781# a_8861_54387# a_10493_52781# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X617 vdd a_7057_34366# a_7257_35054# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=5.16e+06u w=1e+06u l=1e+06u
X618 vdd a_16019_26544# a_15161_31718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X619 a_34723_6373# vss sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=4e+06u
X620 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X621 vdd a_8735_54512# a_9977_51123# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X622 a_43124_15781# vb_3_ a_40013_15426# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X623 vss a_22146_16137# a_22146_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X624 a_7149_30931# a_7257_35054# a_16019_27456# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X625 avdd ibn_0_ a_27033_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X626 a_9215_52237# a_9185_52211# vss vss sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X627 a_21015_51763# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X628 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X629 a_22146_16137# a_21230_16137# a_21230_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X630 a_46648_5440# a_46202_5068# a_46552_5440# vss sky130_fd_pr__nfet_01v8 ad=2.802e+11p pd=2.2e+06u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X631 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X632 a_27549_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X633 a_6416_39560# refsel vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X634 a_14147_17413# a_14605_15614# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X635 a_14147_17185# a_14147_17185# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X636 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X637 vdd a_16019_26544# a_15161_31718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X638 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X639 a_21793_19294# a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X640 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X641 a_40013_15426# a_40013_15754# a_40013_15426# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X642 a_43124_15781# ibp_2_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X643 vdd a_8915_50061# a_9978_51925# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.087e+11p ps=1.36e+06u w=420000u l=150000u
X644 a_16534_48421# a_15795_54391# vb_2_ vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X645 a_21015_51763# a_21015_51763# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X646 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X647 vdd a_14147_17185# a_14147_17413# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X648 a_9091_54413# a_8737_54413# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X649 a_10493_52781# a_10383_52897# a_10533_55475# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X650 a_43124_15781# ibp_2_ vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X651 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X652 a_28184_49195# a_28184_49195# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X653 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X654 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X655 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X656 vdd a_21333_59018# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X657 vss a_8735_54512# a_10533_56019# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X658 a_9185_52211# a_9521_52211# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X659 a_47117_5440# a_46036_5068# a_46770_5036# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.176e+11p pd=1.4e+06u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X660 a_21230_16137# a_21230_16137# a_21230_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X661 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X662 a_11926_4549# a_12242_4494# a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X663 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X664 a_9065_53299# a_9039_52781# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X665 a_21333_59018# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X666 vss a_21272_47107# a_21272_47107# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X667 a_17146_5558# a_18412_7690# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X668 vss a_32117_14563# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X669 a_15338_13967# a_14605_15614# a_14147_17185# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=6.32e+06u w=500000u l=8e+06u
X670 a_14147_17413# a_14147_17185# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X671 vdd a_9506_17973# a_9506_17973# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X672 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X673 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X674 a_8871_56045# tbctl_0_ vss vss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X675 a_7080_26645# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X676 vss a_9975_50061# a_10143_50061# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X677 vss a_21230_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X678 avdd a_9033_7909# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X679 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X680 a_36712_33396# a_37870_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X681 a_39286_5164# a_38936_5164# a_39191_5164# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X682 vss a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X683 vss a_8861_54387# a_9521_52211# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X684 vss ibp_1_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X685 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X686 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X687 a_15161_30727# a_16019_26544# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X688 a_10803_51693# a_8915_50061# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X689 dvdd a_46031_5758# a_46036_5606# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X690 a_16534_48421# a_16071_54391# vb_2_ vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X691 a_46814_5428# a_46770_5036# a_46648_5440# vss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X692 a_47226_5440# a_46036_5068# a_47117_5440# vss sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=1.422e+11p ps=1.51e+06u w=360000u l=150000u
X693 a_21088_54984# a_21088_54984# a_21030_55081# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X694 vdd a_9506_17973# a_8302_16888# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X695 a_21533_59718# a_28184_49195# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X696 a_40013_15754# a_40013_15754# a_40013_15754# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X697 a_8302_16888# a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X698 a_21531_53226# ibp_0_ a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X699 a_21015_51763# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X700 vss a_6880_26619# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X701 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X702 a_9697_51123# a_10435_54957# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X703 a_16534_48421# a_17233_54391# vb_3_ vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X704 a_29267_5405# a_27549_7238# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X705 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X706 a_21015_51763# a_16534_48421# a_21531_53226# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X707 a_8861_54387# a_9065_53299# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X708 vss a_22146_16137# a_22146_17193# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X709 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X710 a_15161_30727# a_16019_26544# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X711 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X712 a_17509_57376# a_17233_57376# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X713 a_22146_17193# a_21230_16137# ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X714 vdd a_21333_59018# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X715 a_21333_59018# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X716 a_9567_53869# a_9697_51123# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X717 vss a_47292_4278# a_47856_3974# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X718 vdd a_10803_51693# a_8735_54512# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X719 a_34011_6373# a_33655_6373# a_29267_5405# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X720 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X721 a_39028_33396# a_37484_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X722 vdd a_8861_54387# a_9473_51399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X723 a_9650_54957# a_9473_54965# vss vss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X724 vss a_40402_5164# a_40757_5164# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X725 ibnbas ibnbas ibnbas vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X726 vss a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X727 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X728 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X729 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X730 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X731 vdd a_9185_52211# a_9215_52237# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X732 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X733 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X734 vdd a_10197_56019# a_10227_56045# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X735 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X736 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X737 a_46340_4145# a_46031_4670# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X738 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X739 vdd a_21030_55081# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X740 vdd a_28184_48339# tbout vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X741 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X742 vbg a_7304_39565# vbg_ext vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X743 a_21088_54984# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X744 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X745 ibnbas ibnbas ibnbas vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X746 a_46031_4670# a_47292_4278# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X747 vdd a_9473_54965# a_9650_54957# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X748 a_28184_49195# a_28184_49195# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X749 vdd a_11221_53325# a_11398_53325# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X750 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X751 a_16534_48421# a_17509_54391# vb_3_ vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X752 vss a_9065_53299# a_8861_54387# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X753 a_28184_49195# ibp_0_ a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X754 vss a_10895_50605# a_11063_50605# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X755 dvdd a_47117_5440# a_47292_5366# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X756 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X757 a_9033_7909# a_9033_7909# a_9033_7909# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X758 a_43124_15781# ibp_2_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X759 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X760 a_9039_52781# a_8871_52781# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X761 a_10493_52781# a_8861_54387# a_10773_52781# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X762 a_40013_15426# a_40013_15754# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X763 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X764 a_8302_16888# a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X765 a_21015_51763# tbout a_21531_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X766 a_8735_54512# a_10803_51693# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X767 a_9215_52237# a_9185_52211# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X768 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X769 a_7080_26645# a_6949_29442# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X770 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X771 vss ibp_2_ ibp_2_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X772 a_21015_51763# a_21015_51763# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X773 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X774 a_7149_30931# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X775 a_21793_19742# a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X776 a_15338_13967# a_14605_15614# a_14147_17185# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X777 a_9697_51123# a_10435_54957# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X778 a_35079_6373# vss sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=4e+06u
X779 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X780 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X781 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X782 a_6633_29468# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X783 vss a_10435_54957# a_9697_51123# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X784 ibp_3_ a_14147_17413# a_21793_20414# vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=3.16e+06u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X785 tbout a_28184_48339# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X786 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X787 a_47756_6694# a_46927_6694# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X788 a_34011_6373# vss sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=4e+06u
X789 a_21257_48618# tbout a_21333_59018# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X790 vss a_6880_26619# a_6880_26619# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X791 a_46340_4731# a_46031_5294# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X792 a_8302_16888# a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X793 a_7257_35054# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X794 a_8915_50061# a_8737_50061# vss vss sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X795 a_47279_4884# a_46202_4518# a_47117_4518# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X796 a_14147_17413# a_14605_15614# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X797 vdd a_10197_55475# a_10227_55501# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X798 a_10533_55475# a_10383_52897# a_10493_52781# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X799 a_40013_15426# a_40013_15426# a_40013_15426# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X800 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X801 vdd a_7057_34366# a_7057_34366# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X802 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X803 a_46031_5294# a_47292_4492# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X804 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X805 a_29435_32656# a_30910_31724# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X806 ibp_2_ ibp_2_ ibp_2_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X807 a_38642_33396# a_37870_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X808 vdd a_9185_52211# a_9215_52237# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X809 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X810 a_14147_17413# a_14605_15614# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X811 vss vdd w_42506_30499# w_42506_30499# sky130_fd_pr__pfet_01v8 ad=4.12764e+14p pd=4.31541e+09u as=0p ps=0u w=1e+06u l=1e+06u
X812 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X813 a_21793_19966# a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X814 a_47267_6832# a_47292_5580# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X815 a_27033_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X816 a_10090_50965# a_9039_52781# a_10018_50965# vss sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=0p ps=0u w=420000u l=150000u
X817 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X818 a_21333_59018# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X819 vss a_9975_50061# a_10143_50061# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X820 vss a_8735_54512# a_9977_51123# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X821 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X822 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X823 a_21531_51763# ibp_0_ a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X824 a_9785_4482# ibp_1_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X825 a_40013_15754# a_40013_15754# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X826 vss a_47292_4492# a_47856_4518# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X827 a_29277_29476# bgtrim_3_ a_30910_30664# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X828 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X829 a_8121_17110# a_8121_17110# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=300000u
X830 a_40013_15426# a_40013_15754# a_40013_15426# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X831 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X832 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X833 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X834 a_9039_52781# a_8871_52781# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X835 dvdd a_47756_6694# clksys dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.12e+12p ps=1.024e+07u w=1e+06u l=150000u
X836 vdd a_10143_50061# a_17233_48421# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X837 a_7149_30931# a_6949_30834# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X838 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X839 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X840 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X841 a_21533_59718# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X842 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X843 a_10533_56019# a_8735_54512# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X844 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X845 a_10383_52897# a_9697_51123# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X846 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X847 vdd a_8735_54512# a_9761_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X848 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X849 vdd a_8933_54387# a_10435_54957# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X850 vss a_6880_26619# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X851 dvdd a_47292_5580# a_47279_5972# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X852 vb_2_ a_32117_17939# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X853 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X854 a_11926_4549# a_11926_4549# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X855 a_47292_4492# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X856 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X857 vss rstn a_39548_5164# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X858 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X859 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X860 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X861 a_7080_26645# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X862 a_9521_52211# a_8861_54387# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X863 a_27549_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X864 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X865 a_16534_48421# a_15795_51406# dvdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X866 vss a_11063_50605# a_15795_51406# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X867 vdd a_9506_17973# a_9506_17973# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X868 vss a_9091_54413# a_9473_54965# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X869 a_21230_16137# a_21230_16137# a_22146_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X870 a_6880_26619# a_7257_35054# a_7257_35054# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X871 a_16196_13967# ibpbas a_15338_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X872 a_22146_16137# a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X873 a_40013_15754# a_40013_15754# a_40013_15754# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X874 a_10227_56045# a_10197_56019# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X875 a_6633_29468# a_6949_30834# a_7149_30931# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X876 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X877 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X878 avdd a_9033_7909# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X879 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X880 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X881 vss vss vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X882 a_39112_16790# a_37846_18922# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X883 vss a_6880_26619# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X884 vss a_46897_6668# a_46927_6694# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X885 a_11398_53325# a_11221_53325# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X886 vss a_9065_53299# a_8861_54387# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X887 a_8871_52781# tbctl_1_ vss vss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X888 vdd a_9506_17973# a_9506_17973# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X889 vdd a_11926_4549# a_11926_4549# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X890 a_16019_27456# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X891 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X892 vdd a_9506_17973# a_8302_16888# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X893 a_28184_49195# a_28184_49195# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X894 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X895 a_29277_29476# bgtrim_9_ a_30910_33844# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X896 a_9185_52211# a_9521_52211# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X897 a_17568_5558# a_17990_7690# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X898 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X899 vdd a_8915_50061# a_10803_51693# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X901 vb_4_ a_32117_17095# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X902 vss vss a_29277_29476# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=0p
X903 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X904 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X905 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X906 a_46660_5062# a_46036_5068# a_46552_5440# dvdd sky130_fd_pr__pfet_01v8_hvt ad=3.402e+11p pd=3.3e+06u as=0p ps=0u w=420000u l=150000u
X907 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X908 a_8302_16888# a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X909 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X910 a_46770_3948# a_46552_4352# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.583e+11p pd=2.37e+06u as=0p ps=0u w=840000u l=150000u
X911 a_8861_54387# a_9065_53299# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X912 a_46457_5606# a_46340_5819# vss vss sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X913 vdd a_10435_54957# a_9697_51123# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X914 vb_3_ a_32117_17939# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X915 a_39028_33396# a_39414_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X916 a_16534_48421# a_17233_51406# vb_4_ vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X917 a_27033_7238# en_clk_int a_33084_7058# avdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X918 a_40757_5164# a_40402_5164# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X919 vdd a_10895_50605# a_11063_50605# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X920 a_9697_51123# a_10435_54957# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X921 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X922 a_46927_6694# a_46897_6668# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X923 vss a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X924 a_21533_59718# a_28184_49195# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X925 a_23557_20190# a_14147_17413# ibp_2_ vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X926 dvdd a_46770_5036# a_46660_5062# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X927 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X928 vss a_21230_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X929 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X930 a_8735_54512# a_10803_51693# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X931 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X932 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X933 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X934 vss a_10197_56019# a_10227_56045# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X935 a_16019_27456# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X936 a_43124_15781# a_37846_16790# a_40013_15754# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X937 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X938 a_16019_27456# ibnbas a_15161_31718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X939 a_10227_55501# a_10197_55475# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X940 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X941 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X942 vdd a_16019_27456# vbg_int vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.45e+12p ps=1.116e+07u w=4e+06u l=1e+06u
X943 vss a_9185_52211# a_9215_52237# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X944 a_6633_29468# a_6949_29442# a_7080_26645# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X945 vdd a_10227_56045# a_17233_57376# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X946 vss a_27549_7238# a_29267_5405# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X947 a_11926_4549# a_12242_4494# a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X948 ibn_0_ a_21230_16137# ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=2.064e+07u as=0p ps=0u w=1e+06u l=2e+06u
X949 a_34367_6373# vss sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=4e+06u
X950 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X951 a_10227_56045# a_10197_56019# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X952 vdd a_21333_59018# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X953 a_9371_53985# a_8861_54387# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X954 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X955 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X956 a_10143_50061# a_9975_50061# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X957 a_43124_15781# a_37846_16790# a_40013_15754# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X958 a_47292_4278# a_47117_4352# a_47471_4340# vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X959 a_16019_26544# ibnbas a_15161_30727# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X960 a_14147_17413# a_14605_15614# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X961 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X962 a_7149_30931# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X963 a_21333_59018# tbout a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X964 a_6880_26619# a_7257_35054# a_7257_35054# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X965 a_21533_59718# a_28184_49195# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X966 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X967 dvdd a_39851_5164# a_40026_5138# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X968 vss a_6880_26619# a_6880_26619# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X969 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X970 a_9785_4482# vb_2_ a_9033_7909# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X971 a_21257_48618# a_16534_48421# a_21533_59718# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X972 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X973 vdd a_9831_50605# a_9931_50721# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X974 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X975 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X976 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X977 a_9183_51693# a_9013_51693# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X978 a_8861_54387# a_9065_53299# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X979 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X980 dvdd a_47292_4492# a_47856_4518# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X981 vdd a_10435_54957# a_9697_51123# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X982 vdd a_21333_59018# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X983 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X984 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X985 a_28184_49195# a_28184_49195# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X986 vss tbctl_0_ a_8871_56045# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X987 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X988 a_10143_50061# a_9975_50061# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X989 vdd a_10895_50605# a_11063_50605# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X990 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X991 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X992 ibp_1_ ibp_1_ ibp_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X993 a_48035_3974# a_47856_3974# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X994 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X995 a_28184_49195# ibp_0_ a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X996 a_9975_50061# a_9650_54957# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X997 dvdd a_38617_5164# a_38770_5164# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X998 dvdd en_clkdiv a_47409_7016# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X999 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1000 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1001 vdd a_11063_50605# a_15795_51406# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1002 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1003 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1004 a_10227_55501# a_10197_55475# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1005 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1006 a_15161_30727# ibnbas a_16019_26544# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1007 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1008 a_46457_5428# a_46340_5233# vss vss sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X1009 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1010 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1011 a_7057_34366# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1012 vdd a_14147_17413# a_14605_15614# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1013 vdd a_14147_17185# a_14147_17413# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X1014 vss a_8871_56045# a_8933_54387# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X1015 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1016 vss a_21272_47107# a_21088_54984# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1017 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1018 a_21257_48618# a_21257_48618# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1019 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1020 dvdd a_47756_6694# clksys dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1021 a_10197_56019# a_10533_56019# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1022 vss en_clkdiv a_47396_6694# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1023 a_15161_31718# ibnbas a_16019_27456# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1024 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1025 avdd a_9033_7909# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1026 a_15161_30727# a_16019_26544# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1027 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1028 vss a_47756_6694# clksys vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1029 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1030 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1031 a_6633_29468# a_6633_29468# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1032 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1033 a_46031_4206# a_46069_6668# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1034 vss a_6880_26619# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1035 a_10143_50061# a_9975_50061# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X1036 vdd a_8871_52781# a_9039_52781# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1037 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1038 a_16071_48421# a_15795_48421# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1039 vss a_9473_54965# a_9650_54957# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1040 vdd a_10073_52389# a_9013_51925# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1041 vdd a_14147_17185# a_14147_17185# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=1e+07u
X1042 vss a_11221_50213# a_11221_50061# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1043 a_15161_30727# a_16019_26544# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1044 dvdd a_39504_5406# a_39394_5530# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1045 a_47292_4492# a_47117_4518# a_47471_4518# vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1046 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1047 vb_5_ a_32117_16251# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1048 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1049 ibpbas ibpbas vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1050 a_46660_4884# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1051 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1052 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1053 a_8861_54387# a_9065_53299# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1054 a_15338_13967# vbg a_14147_17413# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=6.32e+06u w=500000u l=8e+06u
X1055 vdd a_14147_17413# a_23557_19294# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1056 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1057 a_9697_51123# a_10435_54957# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1058 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1059 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1060 a_21533_59718# a_28184_49195# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1061 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1062 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1063 a_40013_15754# a_37846_16790# a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1064 a_21531_53226# ibp_0_ a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1065 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1066 a_29267_5405# a_27549_7238# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1067 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1068 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1069 vss a_27549_7238# a_27549_7238# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1070 vss a_6880_26619# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1071 vss a_21272_47107# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1072 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1073 a_10197_55475# a_10533_55475# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1074 a_46202_5606# a_46036_5606# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1075 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1076 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1077 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1078 vss a_9185_52211# a_9215_52237# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1079 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1080 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1081 vdd a_9506_17973# a_9506_17973# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1082 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1083 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1084 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1085 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1086 a_29435_36896# a_30910_35964# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1087 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1088 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1089 a_40013_15754# a_37846_16790# a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1090 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1091 vss a_6416_39560# a_7028_39565# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1092 a_21015_51763# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1093 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1094 clksys a_47756_6694# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1095 vss a_8933_54387# a_10435_54957# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1096 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1097 a_28184_48339# a_28184_48339# a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1098 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1099 a_28184_49195# a_28184_49195# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1100 vss a_8737_50061# a_8915_50061# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1101 a_21531_51763# ibp_0_ a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1102 tbout a_28184_48339# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X1103 a_10227_56045# a_10197_56019# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1104 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1105 a_38642_33396# a_39800_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1106 vss a_27549_7238# a_27549_7238# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1107 a_33084_7058# en_clk_int a_33084_6373# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1108 vb_5_ a_32117_15407# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1109 vdd a_7057_34366# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1110 a_9785_4482# ibp_1_ vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1111 a_40013_15754# a_37846_16790# a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1112 vdd a_9065_53299# a_8861_54387# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1113 a_9521_52211# a_9977_51123# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1114 vss a_9650_54957# a_9975_50061# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1115 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1116 a_11063_50605# a_10895_50605# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1117 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1118 avdd ibn_0_ a_27549_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1119 a_40186_33396# a_39800_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1120 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1121 a_40026_5138# a_39851_5164# a_40205_5164# vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1122 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1123 avdd ibn_0_ a_27033_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1124 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1125 a_29277_29476# bgtrim_5_ a_30910_31724# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1126 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1127 a_16534_48421# a_15795_48421# vss vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1128 vss a_8933_54387# a_8891_54413# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X1129 a_21533_59718# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1130 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1131 a_46814_4340# a_46770_3948# a_46648_4352# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X1132 a_16019_27456# a_7257_35054# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1133 vss a_8871_56045# a_8933_54387# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1134 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1135 ibn_0_ a_21230_16137# a_23062_15785# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1136 ibp_1_ ibp_1_ ibp_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1137 a_16071_57376# a_15795_57376# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1138 dvdd a_46031_4670# a_46036_4518# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1139 vbg_int a_16019_27456# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1140 a_23062_15785# a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1141 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1142 vdd a_10197_56019# a_10227_56045# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1143 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1144 a_46031_4206# a_46069_6668# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1145 a_46552_4352# a_46202_3980# a_46457_4340# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.449e+11p pd=1.53e+06u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X1146 a_46202_5068# a_46036_5068# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1147 ibpbas ibpbas vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1148 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1149 a_17509_51406# a_17233_51406# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1150 a_21015_51763# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1151 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1152 a_7057_34366# ibnbas ibnbas vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1153 a_29435_32656# a_30910_32784# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1154 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1155 a_21793_20414# a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1156 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1157 avdd a_9033_7909# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1158 vdd a_9975_50061# a_10143_50061# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1159 a_9855_52053# a_8933_54387# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1160 a_29435_32656# bgtrim_6_ a_29277_29476# vss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1161 vss vss a_29277_29476# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=0p
X1162 clksys a_47756_6694# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1163 avdd ibn_0_ a_27549_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1164 a_47117_4518# a_46202_4518# a_46770_4760# vss sky130_fd_pr__nfet_01v8 ad=1.422e+11p pd=1.51e+06u as=0p ps=0u w=360000u l=150000u
X1165 a_21230_16137# a_21230_16137# a_21230_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1166 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1167 a_21257_48618# a_16534_48421# a_21533_59718# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1168 a_14147_17413# vbg a_15338_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X1169 vss vss vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1170 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1171 vdd a_14147_17413# a_23557_19742# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1172 a_21531_51763# tbout a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1173 a_7057_34366# ibnbas ibnbas vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1174 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1175 avdd ibn_0_ ibn_0_ avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1176 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1177 vdd a_9065_53299# a_8861_54387# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1178 a_28184_48339# a_28184_48339# a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1179 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1180 a_9697_51123# a_10435_54957# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1181 a_16534_48421# a_17233_48421# vbg vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1182 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1183 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1184 vss tbctl_1_ a_8871_52781# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1185 a_9033_7909# vb_2_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1186 a_46031_4670# a_47292_4278# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1187 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1188 vss ibpbas ibpbas vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1189 vdd a_21030_55081# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1190 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1191 a_40581_5164# a_40026_5138# vss vss sky130_fd_pr__nfet_01v8 ad=2.015e+11p pd=1.92e+06u as=0p ps=0u w=650000u l=150000u
X1192 vdd a_10197_55475# a_10227_55501# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1193 a_46202_5606# a_46036_5606# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1194 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1195 a_28184_49195# a_28184_49195# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1196 a_7149_30931# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1197 vss a_40445_30630# a_16019_27456# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1198 ibp_0_ ibp_0_ a_21272_47107# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1199 a_46770_5036# a_46552_5440# vss vss sky130_fd_pr__nfet_01v8 ad=1.998e+11p pd=1.97e+06u as=0p ps=0u w=640000u l=150000u
X1200 vdd a_14147_17413# a_23557_19966# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1201 a_29277_29476# bgtrim_11_ a_30910_34904# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1202 vss a_40026_5138# a_40581_5164# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1203 vss a_8871_52781# a_9039_52781# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1204 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1205 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1206 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1207 a_48035_4518# a_47856_4518# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1208 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1209 avdd a_9033_7909# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1210 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1211 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1212 vss a_10435_54957# a_9697_51123# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1213 a_16019_26544# a_7257_35054# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1214 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1215 a_27549_7238# a_27549_7238# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1216 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1217 vb_0_ a_32117_19627# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1218 a_15161_31718# ibnbas a_16019_27456# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1219 a_46814_4518# a_46770_4760# a_46648_4518# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.802e+11p ps=2.2e+06u w=420000u l=150000u
X1220 ibn_0_ a_21230_16137# ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1221 a_21257_48618# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1222 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1223 vdd a_9975_50061# a_10143_50061# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1224 a_9785_4482# vb_2_ a_9033_7909# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1225 a_27033_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1226 a_9705_51925# a_9978_51925# a_9936_52053# vss sky130_fd_pr__nfet_01v8 ad=1.07825e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1227 a_10227_56045# a_10197_56019# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1228 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1229 vss a_8861_54387# a_10533_56019# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1230 vss vss vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1231 a_9785_4482# vb_2_ a_9033_7909# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1232 a_17568_5558# a_16302_7690# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1233 a_10533_56019# a_9697_51123# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1234 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1235 a_47279_5062# a_46202_5068# a_47117_5440# dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1236 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1237 a_43124_15781# vb_3_ a_40013_15426# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1238 a_15161_30727# ibnbas a_16019_26544# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1239 a_29435_35836# bgtrim_12_ a_29277_29476# vss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1240 a_46568_6694# clkext a_46069_6668# vss sky130_fd_pr__nfet_01v8 ad=1.155e+11p pd=1.39e+06u as=3.465e+11p ps=2.49e+06u w=420000u l=150000u
X1241 a_46648_4352# a_46202_3980# a_46552_4352# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X1242 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1243 a_46552_5440# a_46036_5068# a_46457_5428# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1244 a_7080_26645# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1245 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1246 vdd a_8933_54387# a_8737_54413# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X1247 a_29435_29476# a_30910_29604# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1248 clksys a_47756_6694# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1249 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1250 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1251 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1252 a_28184_48339# a_28184_48339# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1253 a_28184_48339# ibp_0_ a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1254 a_21088_54984# a_21088_54984# a_21030_55081# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1255 dvdd a_40013_15426# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1256 a_21015_51763# tbout a_21531_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1257 a_14147_17413# vbg a_15338_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X1258 a_29435_35836# a_30910_34904# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1259 vss a_10227_55501# a_15795_57376# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1260 vdd a_21333_59018# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1261 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1262 a_8742_39565# a_8466_39565# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1263 vb_1_ a_32117_19627# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1264 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1265 a_17509_51406# a_17233_51406# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1266 a_27549_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1267 a_21230_16137# a_14147_17413# a_21793_19518# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1268 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1269 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1270 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1271 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1272 dvdd a_47292_4492# a_47279_4884# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1273 a_28184_48339# a_28184_48339# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1274 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1275 a_47292_5366# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1276 vdd a_9975_50061# a_10143_50061# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1277 a_39074_5377# a_40581_5164# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1278 a_46457_4340# a_46340_4145# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1279 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1280 vdd a_21030_55081# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1281 a_39960_5164# a_38770_5164# a_39851_5164# vss sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X1282 vdd a_9013_51925# a_9013_51693# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X1283 dvdd a_47292_5366# a_47856_5062# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1284 a_40013_15754# a_40013_15754# a_40013_15754# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1285 clksys a_47756_6694# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1286 a_47075_6846# en_clkdiv vss vss sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X1287 a_8933_54387# a_8871_56045# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1288 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1289 a_8871_52781# tbctl_1_ vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1290 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1291 a_40572_33396# a_39414_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1292 vss ibp_1_ ibp_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1293 w_42506_30499# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1294 a_8737_54413# a_8861_54387# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1295 a_47226_4352# a_46036_3980# a_47117_4352# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1296 ibp_2_ ibp_2_ vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1297 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1298 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1299 ibp_0_ ibp_0_ a_21272_47107# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1300 vdd a_8915_50061# a_9931_50721# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1301 a_10803_51693# a_8915_50061# vss vss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X1302 a_9831_50605# a_8933_54387# vss vss sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1303 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1304 vss a_39534_18922# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1305 a_7149_30931# a_6949_30834# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1306 vss a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1307 a_11926_4549# a_11926_4549# a_11926_4549# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1308 a_46648_5606# a_46202_5606# a_46552_5606# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.188e+11p ps=1.38e+06u w=360000u l=150000u
X1309 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1310 vss a_11221_50061# a_11398_50061# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1311 dvdd a_40013_15426# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1312 a_21333_59018# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1313 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1314 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1315 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1316 a_21272_47107# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1317 vss a_9705_51925# a_9105_50837# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1318 vss a_8871_52781# a_9039_52781# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1319 avdd ibn_0_ a_27549_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1320 w_42506_30499# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1321 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1322 a_7080_26645# a_6949_29442# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1323 a_8915_50061# a_8737_50061# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1324 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1325 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1326 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1327 a_6633_29468# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1328 vss a_10435_54957# a_9697_51123# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1329 vss a_9039_52781# a_10346_52217# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.0785e+11p ps=1.36e+06u w=420000u l=150000u
X1330 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1331 a_29435_31596# a_30910_31724# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1332 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1333 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1334 a_39394_5530# a_38770_5164# a_39286_5164# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1335 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1336 a_10197_56019# a_10533_56019# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1337 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1338 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1339 vss ibpbas a_16196_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1340 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1341 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1342 a_9033_7909# a_11926_4549# a_9033_7909# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1343 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1344 vss a_9215_52237# a_17233_51406# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1345 a_28184_48339# ibp_0_ a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1346 a_7149_30931# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1347 ibp_2_ ibp_2_ ibp_2_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1348 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1349 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1350 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1351 avdd a_16724_7690# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1352 vbg a_8466_39565# vbg_int vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1353 a_9033_7909# a_9033_7909# a_9033_7909# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1354 a_29435_29476# a_29277_29476# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1355 a_46552_5606# a_46202_5606# a_46457_5606# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X1356 a_27549_7238# a_27549_7238# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1357 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1358 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1359 a_21333_59018# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1360 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1361 a_47226_5606# a_46036_5606# a_47117_5606# vss sky130_fd_pr__nfet_01v8 ad=1.338e+11p pd=1.5e+06u as=0p ps=0u w=360000u l=150000u
X1362 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1363 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1364 avdd ibn_0_ a_27033_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1365 dvdd a_40013_15426# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1366 vdd a_11926_4549# a_11926_4549# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1367 a_11221_50213# a_11129_51149# vss vss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1368 a_16019_26544# a_7257_35054# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1369 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1370 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1371 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1372 vss a_22146_16137# a_22146_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1373 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1374 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1375 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1376 a_22146_16137# a_21230_16137# a_21230_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1377 vss a_47756_6694# clksys vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1378 vdd a_8121_17110# a_8302_16888# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=300000u
X1379 dvdd a_40402_5164# a_40757_5164# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1380 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1381 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1382 dvdd a_46897_6668# a_46927_6694# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1383 a_46031_5294# a_47292_4492# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1384 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1385 a_9761_53869# a_9697_51123# a_9481_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X1386 a_15338_13967# vbg a_14147_17413# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X1387 a_23557_19294# a_14147_17413# ibp_1_ vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1388 a_10435_54957# a_8933_54387# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1389 a_43124_15781# ibp_2_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1390 a_8891_54413# a_8861_54387# a_8819_54413# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1391 vss a_9275_50605# a_11221_53325# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1392 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1393 a_11063_50605# a_10895_50605# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1394 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1395 vss a_10287_50605# a_11129_51149# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X1396 vss ibp_2_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1397 a_40186_33396# a_41344_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1398 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1399 ibn_0_ a_21230_16137# a_23062_16841# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1400 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1401 a_46457_4340# a_46340_4145# vss vss sky130_fd_pr__nfet_01v8 ad=1.32e+11p pd=1.49e+06u as=0p ps=0u w=420000u l=150000u
X1402 a_23062_16841# a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1403 a_10143_50061# a_9975_50061# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1404 a_39053_30692# a_16019_27456# vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1405 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1406 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1407 a_39074_5377# a_40581_5164# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1408 a_6633_29468# a_6949_29442# a_7080_26645# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1409 a_7080_26645# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1410 vdd a_10283_54413# a_15795_54391# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1411 a_27549_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1412 vss a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1413 vdd a_9705_51925# a_9105_50837# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1414 ibp_1_ ibp_1_ ibp_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1415 ibp_1_ ibp_1_ vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1416 a_21531_51763# tbout a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1417 a_8933_54387# a_8871_56045# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1418 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1419 vss a_6880_26619# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1420 clksys a_47756_6694# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1421 ibn_0_ a_21230_16137# ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1422 a_28184_49195# a_28184_49195# a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1423 a_21333_59018# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1424 vdd a_8735_54512# a_8737_54413# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1425 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1426 a_11926_4549# a_12242_4494# a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1427 vdd a_7057_34366# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1428 dvdd a_47292_5580# a_47856_5606# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1429 a_16196_13967# ibpbas vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1430 vdd en_ldo_dig a_47886_16107# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1431 a_8735_54512# a_10803_51693# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1432 a_9481_53869# a_9371_53985# a_9567_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X1433 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1434 a_34367_6373# a_34011_6373# a_27033_7238# avdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1435 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1436 a_21257_48618# a_21257_48618# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1437 dvdd a_40026_5138# a_40581_5164# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1438 a_46069_6668# a_40581_5164# a_46278_6694# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1439 vdd a_7057_34366# a_7257_35054# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1440 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1441 vss vss vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1442 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1443 a_43124_15781# vb_3_ a_40013_15426# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1444 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1445 a_21030_55081# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1446 a_9039_52781# a_8871_52781# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1447 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1448 a_40013_15754# a_37846_16790# a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1449 a_15338_13967# ibpbas a_16196_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1450 vb_3_ a_32117_17095# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1451 a_33004_6347# vss sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=4e+06u
X1452 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1453 clksys a_47756_6694# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1454 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1455 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1456 a_9975_50061# a_9650_54957# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1457 a_29435_31596# a_30910_30664# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1458 a_6949_30834# a_34396_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1459 a_10223_52243# a_8915_50061# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1460 a_10435_54957# a_8933_54387# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1461 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1462 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1463 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1464 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1465 a_21531_53226# a_16534_48421# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1466 a_9785_4482# a_12242_4494# a_11926_4549# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1467 a_46660_5062# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1468 a_6633_29468# a_6633_29468# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1469 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1470 a_16019_27456# a_7257_35054# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1471 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1472 a_11063_50605# a_10895_50605# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1473 a_14147_17413# a_14605_15614# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1474 a_6633_29468# a_6949_30834# a_7149_30931# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1475 a_21531_53226# a_16534_48421# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1476 a_27549_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1477 a_46770_5848# a_46552_5606# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1478 vss a_40026_5138# a_40402_5164# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1479 vdd a_21333_59018# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1480 a_21333_59018# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1481 a_40757_5164# a_40402_5164# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1482 vdd a_9215_52237# a_17233_51406# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1483 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1484 a_11398_50061# a_11221_50061# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1485 a_40026_5138# rstn dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1486 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1487 avdd ibn_0_ a_27549_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1488 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1489 vdd tbctl_1_ a_8871_52781# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1490 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1491 vss a_21230_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1492 a_9039_52781# a_8871_52781# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1493 a_37082_4920# a_33004_6347# avdd avdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1494 dvdd a_46069_6668# a_46031_4206# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1495 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1496 a_46457_4518# a_46340_4731# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1497 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1498 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1499 a_43124_15781# ibp_2_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1500 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1501 a_9506_17973# a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1502 vss a_10197_56019# a_10227_56045# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1503 vdd a_14147_17413# a_14605_15614# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1504 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1505 a_46457_5606# a_46340_5819# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1506 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1507 a_10283_54413# a_10117_54413# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=5.4e+11p pd=5.08e+06u as=0p ps=0u w=1e+06u l=150000u
X1508 vss a_9697_51123# a_10533_56019# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1509 a_39053_30692# a_40958_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1510 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1511 a_7149_30931# a_7257_35054# a_16019_27456# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1512 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1513 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1514 vss a_47756_6694# clksys vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1515 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1516 a_14147_17185# a_14605_15614# a_15338_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X1517 a_6633_29468# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1518 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1519 avdd ibn_0_ a_27033_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1520 a_23557_19742# a_14147_17413# ibp_0_ vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1521 a_28184_48339# a_28184_49195# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1522 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1523 ibnbas ibnbas a_7057_34366# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1524 a_27033_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1525 vdd a_8737_50061# a_8915_50061# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1526 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1527 a_9481_53869# a_9697_51123# a_9761_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1528 vdd a_21333_59018# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1529 vdd a_14147_17413# a_23557_20414# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=3.16e+06u w=500000u l=2e+06u
X1530 vdd a_16019_26544# a_15161_31718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1531 a_29435_36896# bgtrim_14_ a_29277_29476# vss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1532 vdd a_21333_59018# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1533 a_10287_50605# a_9931_50721# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1534 a_8302_16888# a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1535 tbout a_28184_48339# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X1536 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1537 a_46340_5233# a_46031_5758# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1538 ibnbas ibnbas a_7057_34366# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1539 a_10073_52389# a_8915_50061# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1540 a_17509_57376# a_17233_57376# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1541 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1542 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1543 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1544 a_29435_29476# bgtrim_0_ a_29277_29476# vss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1545 a_16071_51406# a_15795_51406# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1546 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1547 a_7149_30931# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1548 vdd a_16019_26544# a_15161_31718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1549 vdd a_21030_55081# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1550 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1551 a_23557_19966# a_14147_17413# ibp_0_ vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1552 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1553 vdd a_9275_50605# a_11221_53325# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1554 vss a_27549_7238# a_29267_5405# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1555 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1556 vss a_21272_47107# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1557 a_28184_49195# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1558 a_46202_3980# a_46036_3980# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1559 a_6416_39560# refsel vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1560 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1561 a_47117_4352# a_46036_3980# a_46770_3948# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1562 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1563 vss a_10197_55475# a_10227_55501# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1564 a_9567_53869# a_9371_53985# a_9481_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1565 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1566 a_21531_53226# ibp_0_ a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1567 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1568 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1569 a_9705_51925# a_9978_51925# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1570 vdd a_21333_59018# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1571 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1572 a_21015_51763# tbout a_21531_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1573 a_35168_33396# a_34782_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1574 a_16019_27456# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1575 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1576 a_27033_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1577 a_10895_50605# a_9183_51693# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X1578 a_21015_51763# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1579 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1580 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1581 a_21533_59718# a_28184_49195# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1582 a_10283_54413# a_10117_54413# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1583 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1584 a_40013_15426# vb_3_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1585 vbg_int a_41344_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1586 a_6633_29468# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1587 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1588 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1589 vss a_6880_26619# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1590 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1591 a_21257_48618# tbout a_21333_59018# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1592 dvdd a_40026_5138# a_40402_5164# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1593 a_11926_4549# a_11926_4549# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1594 vss a_8915_50061# a_10803_51693# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1595 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1596 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1597 vdd a_10895_50605# a_11063_50605# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1598 a_7080_26645# a_7257_35054# a_16019_26544# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1599 a_6633_29468# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1600 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1601 a_7257_35054# a_7257_35054# a_7257_35054# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1602 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1603 a_29435_35836# a_30910_35964# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1604 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1605 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X1606 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1607 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1608 vss vss a_29277_29476# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=0p
X1609 a_47106_6694# a_47075_6846# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1610 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1611 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1612 a_46202_4518# a_46036_4518# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=0p ps=0u w=640000u l=150000u
X1613 vss en_ldo_dig a_47886_16107# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1614 a_34367_6373# a_34011_6373# a_29267_5405# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1615 a_14147_17413# a_14605_15614# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1616 a_48035_5062# a_47856_5062# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1617 a_9039_52781# a_8871_52781# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1618 vss vss vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1619 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1620 vss vss a_29277_29476# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=0p
X1621 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1622 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1623 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1624 a_6633_29468# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1625 ibn_0_ ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1626 a_9697_51123# a_10435_54957# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1627 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1628 a_21015_51763# a_21015_51763# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1629 a_46069_6668# clkext a_46296_7016# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=4.576e+11p ps=2.71e+06u w=640000u l=150000u
X1630 clksys a_47756_6694# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1631 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1632 a_46927_6694# a_46897_6668# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1633 a_21793_19518# a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1634 vss a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1635 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1636 vss a_46927_6694# a_47756_6694# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.176e+11p ps=1.4e+06u w=420000u l=150000u
X1637 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1638 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1639 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1640 a_38690_16790# a_38268_18922# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1641 a_7149_30931# a_6949_30834# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1642 a_27033_7238# ibn_0_ avdd avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1643 vb_6_ a_32117_15407# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1644 a_14605_15614# a_32117_20471# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1645 a_21015_51763# tbout a_21531_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1646 a_21533_59718# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1647 vss a_10383_52897# a_10533_55475# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1648 vdd a_7057_34366# a_7057_34366# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1649 a_10865_53869# a_8735_54512# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1650 a_28184_49195# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1651 a_6949_29442# a_34782_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1652 dvdd a_47117_4352# a_47292_4278# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1653 vss a_21272_47107# a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1654 a_21088_54984# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1655 a_28184_49195# a_28184_49195# a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1656 vdd a_9567_53869# a_10117_54413# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X1657 a_46202_4518# a_46036_4518# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1658 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1659 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1660 tbout a_28184_48339# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X1661 a_21531_53226# ibp_0_ a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1662 a_21531_53226# ibp_0_ a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1663 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X1664 vss a_22146_16137# a_22146_15785# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1665 a_21030_55081# a_21088_54984# a_21088_54984# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1666 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1667 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1668 a_9033_7909# vb_2_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1669 a_22146_15785# a_21230_16137# ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1670 a_29435_30536# a_30910_29604# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1671 vss a_6880_26619# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1672 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1673 vdd w_42506_30499# a_40445_30630# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1674 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1675 a_40445_30630# vbg_int vss vss sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X1676 a_16019_26544# a_16019_26544# a_16019_26544# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1677 a_29267_5405# a_27549_7238# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1678 a_37082_4920# a_33004_6347# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1679 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1680 ibp_1_ a_9033_6762# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=400000u
X1681 a_16071_51406# a_15795_51406# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1682 a_39112_16790# a_39534_18922# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1683 a_7909_13748# vdd vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1684 vss vss a_29277_29476# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=0p
X1685 vss a_21230_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1686 a_9183_51693# a_9013_51693# vss vss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1687 vdd a_8871_56045# a_8933_54387# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1688 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1689 ibn_1_ a_21230_16137# ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1690 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1691 a_40013_15754# a_40013_15754# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1692 vss a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1693 a_16019_26544# a_16019_26544# a_16019_26544# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1694 a_10773_52781# a_8735_54512# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1695 a_7257_35054# a_7257_35054# a_7257_35054# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1696 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1697 vss a_11221_53325# a_11398_53325# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X1698 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1699 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1700 a_47756_6694# a_46927_6694# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1701 a_28184_49195# ibp_0_ a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1702 a_17509_54391# a_17233_54391# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1703 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1704 a_9761_53869# a_8735_54512# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1705 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1706 a_21257_48618# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1707 vdd a_9039_52781# a_9705_51925# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1708 ibn_0_ a_21230_16137# ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1709 a_21257_48618# tbout a_21333_59018# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1710 ibpbas ibpbas vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1711 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1712 ibp_1_ ibp_1_ vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1713 a_10143_50061# a_9975_50061# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1714 dvdd a_47292_5366# a_47279_5062# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1715 a_33655_6373# a_33084_7058# a_27033_7238# avdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1716 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1717 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1718 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1719 dvdd a_47756_6694# clksys dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1720 vdd a_10117_54413# a_10283_54413# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1721 a_9506_17973# a_9506_17973# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1722 vss a_6880_26619# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1723 vss a_8871_56045# a_8933_54387# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1724 vdd a_28184_48339# tbout vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X1725 a_16019_27456# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1726 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1727 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1728 vss a_38617_5164# a_38770_5164# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1729 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1730 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1731 a_7149_30931# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1732 vdd a_21030_55081# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1733 vss a_21272_47107# a_21272_47107# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1734 vss a_47292_5580# a_47226_5606# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1735 a_10227_55501# a_10197_55475# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1736 vss a_11398_50061# a_15795_48421# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1737 a_28184_49195# ibp_0_ a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1738 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1739 a_16534_48421# a_16071_48421# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1740 a_40013_15426# a_40013_15754# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1741 a_7080_26645# a_7257_35054# a_16019_26544# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1742 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1743 vss a_9371_53985# a_9567_53869# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1744 a_6633_29468# a_6949_29442# a_7080_26645# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1745 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1746 vss ibpbas ibpbas vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=4e+06u
X1747 a_10895_50605# a_9183_51693# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1748 vss a_10803_51693# a_8735_54512# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1749 a_38617_5164# a_37082_4920# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1750 a_28184_48339# a_28184_49195# a_21533_59718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1751 vdd a_8871_56045# a_8933_54387# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1752 a_43124_15781# a_37846_16790# a_40013_15754# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1753 w_42506_30499# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1754 a_16019_26544# a_16019_26544# a_16019_26544# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1755 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1756 a_21531_51763# ibp_0_ a_28184_49195# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1757 ibnbas a_8302_16888# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1758 a_35554_33396# a_34396_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1759 ibp_1_ ibp_1_ ibp_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1760 vss a_10227_56045# a_17233_57376# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1761 a_21533_59718# a_28184_49195# a_28184_48339# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1762 a_11926_4549# a_11926_4549# a_11926_4549# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1763 a_46340_5819# a_47267_6832# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1764 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1765 a_47471_5606# rstn vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1766 a_12242_4494# a_18412_7690# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1767 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1768 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1769 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1770 a_16019_26544# a_16019_26544# a_16019_26544# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1771 vss a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1772 vdd a_9183_51693# a_10895_50605# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1773 vdd a_8735_54512# a_10865_53869# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1774 a_10283_54413# a_10117_54413# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1775 vdd a_10117_54413# a_10283_54413# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1776 vss rstn a_46814_5606# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1777 a_21015_51763# a_21015_51763# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1778 a_46770_3948# a_46552_4352# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1779 a_16019_26544# ibnbas a_15161_30727# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1780 avdd ibn_0_ a_27033_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1781 ibp_2_ a_14147_17413# a_21793_20190# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1782 a_46247_6846# clksel dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=1.728e+11p pd=1.82e+06u as=0p ps=0u w=640000u l=150000u
X1783 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1784 a_16534_48421# a_17509_48421# vbg vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1785 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1786 a_46660_3974# a_46036_3980# a_46552_4352# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1787 a_21531_51763# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1788 a_47117_5606# a_46036_5606# a_46770_5848# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.583e+11p ps=2.37e+06u w=420000u l=150000u
X1789 vdd a_40013_15754# a_40013_15426# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1790 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1791 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1792 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1793 a_46552_4518# a_46202_4518# a_46457_4518# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.302e+11p ps=1.46e+06u w=420000u l=150000u
X1794 a_29435_34776# a_30910_34904# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1795 vss a_8735_54512# a_9567_53869# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1796 a_46770_5848# a_46552_5606# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1797 a_16019_27456# ibnbas a_15161_31718# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1798 vss a_46031_5758# a_46036_5606# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1799 dvdd a_46770_3948# a_46660_3974# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1800 a_10533_55475# a_10383_52897# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1801 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1802 a_21333_59018# tbout a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1803 vb_1_ a_32117_18783# vss sky130_fd_pr__res_xhigh_po w=690000u l=2.58e+07u
X1804 a_40013_15426# a_40013_15426# a_40013_15426# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1805 dvdd a_39956_18922# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1806 a_37846_16790# a_38268_18922# vss sky130_fd_pr__res_xhigh_po w=350000u l=8.5e+06u
X1807 vss a_47292_5366# a_47226_5440# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1808 a_21333_59018# a_28184_49195# a_28184_49195# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1809 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1810 vss clksel a_46568_6694# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1811 a_7080_26645# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1812 a_28184_49195# ibp_0_ a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1813 vss a_8915_50061# a_9978_51925# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.0785e+11p ps=1.36e+06u w=420000u l=150000u
X1814 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1815 a_9931_50721# a_9039_52781# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1816 a_7149_30931# a_7257_35054# a_16019_27456# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1817 vdd a_9033_7909# avdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1818 vss a_6880_26619# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1819 a_46552_4352# a_46036_3980# a_46457_4340# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1820 vss a_8915_50061# a_10090_50965# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1821 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1822 a_28184_49195# ibp_0_ a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1823 a_46340_5233# a_46031_5758# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1824 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1825 dvdd a_40013_15426# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1826 vdd a_9650_54957# a_9975_50061# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1827 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1828 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1829 a_39191_5164# a_39074_5377# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1830 a_8933_54387# a_8871_56045# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1831 a_46031_5758# a_47292_5366# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=0p ps=0u w=1e+06u l=150000u
X1832 dvdd a_47756_6694# clksys dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1833 vdd a_40013_15754# a_40013_15754# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1834 a_47471_5428# rstn vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1835 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1836 a_9275_50605# a_9105_50605# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X1837 a_9033_7909# a_11926_4549# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1838 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1839 dvdd a_40013_15426# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1840 a_10227_55501# a_10197_55475# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1841 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1842 a_11398_53325# a_11221_53325# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1843 a_7304_39565# a_7028_39565# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1844 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1845 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1846 a_21333_59018# tbout a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1847 vss rstn a_46814_5428# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1848 vss a_10283_54413# a_15795_54391# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1849 a_35168_33396# a_36326_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1850 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1851 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1852 a_7149_30931# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1853 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1854 vss a_10803_51693# a_8735_54512# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1855 a_38617_5164# a_37082_4920# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X1856 dvdd a_47117_5606# a_47292_5580# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1857 a_47117_5440# a_46202_5068# a_46770_5036# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1858 ibn_1_ a_21230_16137# a_23062_15433# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1859 a_8933_54387# a_8871_56045# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1860 vss vss a_29277_29476# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=0p
X1861 a_14147_17185# a_14605_15614# a_15338_13967# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=8e+06u
X1862 a_23062_15433# a_22146_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1863 vss a_6880_26619# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1864 a_6633_29468# a_6633_29468# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1865 a_21030_55081# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1866 vdd a_11926_4549# a_9033_7909# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1867 a_21531_53226# a_21272_47107# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1868 a_15161_31718# a_16019_26544# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1869 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1870 vss a_46031_5294# a_46036_5068# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1871 a_21015_51763# a_16534_48421# a_21531_53226# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1872 a_33655_6373# a_33084_7058# a_29267_5405# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1873 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1874 vss a_27549_7238# a_29267_5405# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1875 a_9473_51399# a_9697_51123# a_9727_51399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1876 tbout a_28184_48339# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=4e+06u
X1877 a_23557_20414# a_14147_17413# ibp_3_ vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1878 a_21230_16137# a_21230_16137# a_21230_16137# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1879 vdd refsel a_8466_39565# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1880 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1881 a_43124_15781# ibp_2_ vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1882 a_28184_48339# a_28184_48339# a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1883 a_10283_54413# a_10117_54413# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1884 a_46648_4518# a_46202_4518# a_46552_4518# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1885 a_9567_53869# a_9371_53985# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1886 a_15161_31718# a_16019_26544# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1887 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1888 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1889 vdd a_11398_53325# a_17233_54391# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=400000u
X1890 dvdd vss dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1891 a_46552_5606# a_46036_5606# a_46457_5606# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1892 a_21533_59718# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1893 dvdd a_40026_5138# a_40013_5530# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.134e+11p ps=1.38e+06u w=420000u l=150000u
X1894 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1895 vss a_8871_52781# a_9039_52781# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1896 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1897 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1898 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1899 a_16019_27456# a_7257_35054# a_7149_30931# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1900 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1901 vdd a_9039_52781# a_10346_52217# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.087e+11p ps=1.36e+06u w=420000u l=150000u
X1902 a_40013_5530# a_38936_5164# a_39851_5164# dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1903 a_28184_49195# ibp_0_ a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1904 a_28184_49195# ibp_0_ a_21531_51763# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1905 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1906 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1907 a_29435_34776# a_30910_33844# vss sky130_fd_pr__res_high_po w=1.41e+06u l=2.8e+06u
X1908 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1909 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1910 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1911 a_28184_49195# a_28184_49195# a_21333_59018# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1912 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1913 vss dvdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1914 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1915 vss a_22146_16137# a_22146_16841# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1916 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1917 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1918 a_9033_7909# vb_2_ a_9785_4482# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1919 a_22146_16841# a_21230_16137# ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1920 avdd a_9033_7909# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1921 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1922 a_35554_33396# a_35940_36428# vss sky130_fd_pr__res_xhigh_po w=690000u l=1.3e+07u
X1923 a_7080_26645# a_6949_29442# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1924 vss vss a_29277_29476# vss sky130_fd_pr__pnp_05v5_W0p68L0p68 area=0p
X1925 vss a_40026_5138# a_39960_5164# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1926 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X1927 vss a_9567_53869# a_10117_54413# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1928 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1929 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X1930 vss a_10073_52389# a_9013_51925# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X1931 a_46457_4518# a_46340_4731# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1932 a_8933_54387# a_8871_56045# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1933 a_9785_4482# a_12242_4494# a_11926_4549# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1934 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1935 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1936 avdd ibn_0_ a_27033_7238# avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1937 a_46296_7016# a_46247_6846# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1938 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1939 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1940 a_9275_50605# a_9105_50605# vss vss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X1941 vss a_21272_47107# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1942 a_16071_57376# a_15795_57376# vss vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1943 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1944 vdd a_11221_50213# a_11221_50061# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1945 a_29435_30536# bgtrim_2_ a_29277_29476# vss sky130_fd_pr__nfet_01v8 ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=500000u
X1946 a_39191_5164# a_39074_5377# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1947 a_9340_13770# a_9448_14814# vss sky130_fd_pr__res_xhigh_po w=350000u l=7e+06u
X1948 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1949 a_7257_35054# a_7057_34366# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1950 a_9831_50605# a_8933_54387# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1951 a_21533_59718# a_21333_59018# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1952 a_47226_4518# a_46036_4518# a_47117_4518# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1953 a_9506_17973# a_8302_16888# a_9448_14814# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X1954 vss vss vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1955 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1956 a_21257_48618# a_21257_48618# a_21257_48618# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1957 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1958 a_40013_15426# vb_3_ a_43124_15781# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1959 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1960 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1961 a_33084_7058# a_33004_6347# a_27033_7238# avdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=400000u
X1962 a_33004_6347# a_35079_6373# a_27033_7238# avdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=400000u
X1963 vdd a_14147_17413# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
X1964 vss a_21272_47107# a_21531_53226# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1965 vdd a_40013_15426# dvdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1966 vss a_21230_16137# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1967 vss a_6880_26619# a_7080_26645# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1968 vdd a_7057_34366# a_6633_29468# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1969 ibn_1_ a_21230_16137# ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1970 a_10197_55475# a_10533_55475# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X1971 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X1972 dvdd a_40013_15426# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
X1973 a_28184_48339# a_28184_48339# a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1974 a_21531_53226# ibp_0_ a_28184_48339# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=4e+06u
X1975 a_9521_52211# a_9977_51123# a_9727_51399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1976 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1977 a_21015_51763# a_21030_55081# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1978 a_16019_27456# vss sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
X1979 vdd a_21030_55081# a_21015_51763# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1980 a_7080_26645# a_6880_26619# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1981 avdd a_9033_7909# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=500000u
X1982 a_29277_29476# bgtrim_7_ a_30910_32784# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=500000u
X1983 avdd ibn_0_ ibn_0_ avdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1984 a_46770_5036# a_46552_5440# dvdd dvdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1985 a_38936_5164# a_38770_5164# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X1986 vdd a_14147_17413# a_14605_15614# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=500000u l=2e+06u
.ends

