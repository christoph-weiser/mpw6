* SPICE3 file created from decoder3to8.ext - technology: sky130A


* Top level circuit decoder3to8

.subckt decoder3to8 out5 vdd vss out4 out3 out2 out1 out0 out6 out7 in0 in1 in2
X0 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=3.30922e+13p pd=3.6296e+08u as=0p ps=0u w=550000u l=590000u
X1 vdd a_1731_2919# a_671_2455# vdd sky130_fd_pr__pfet_01v8_hvt ad=4.72991e+13p pd=4.6549e+08u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X2 a_1308_5487# a_1131_5495# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_1363_2455# a_1636_2455# a_1594_2583# vss sky130_fd_pr__nfet_01v8 ad=1.07825e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X4 a_841_2223# a_671_2223# vss vss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X5 vdd a_1775_4943# out2 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X6 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X7 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X8 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X9 a_393_5042# a_2461_2223# vss vss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X10 out7 a_1633_591# vss vss sky130_fd_pr__nfet_01v8 ad=5.265e+11p pd=5.52e+06u as=0p ps=0u w=650000u l=150000u
X11 a_477_4943# a_393_5042# a_395_4943# vss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X12 a_1489_1135# a_591_4917# vss vss sky130_fd_pr__nfet_01v8 ad=1.0785e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X13 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X14 vdd a_529_6575# a_591_4917# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X15 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X16 vdd a_591_4917# a_395_4943# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.415e+11p ps=2.83e+06u w=420000u l=150000u
X17 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X18 a_1029_4515# a_519_4917# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X19 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X20 vdd a_1489_1135# a_1589_1251# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X21 vss a_1731_2919# a_671_2455# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X22 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X23 vdd a_529_6575# a_591_4917# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X25 a_1385_1929# a_1635_1653# a_1179_2741# vdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X26 vdd a_393_5042# a_1419_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X27 vdd in0 a_529_6575# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X28 out2 a_1775_4943# vss vss sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X29 a_1355_1653# a_2093_5487# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X30 vdd a_2879_591# out6 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X31 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X32 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X33 vss a_1355_1653# a_1225_4399# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X34 a_1748_1495# a_697_3311# a_1676_1495# vss sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X35 a_1139_4399# a_1355_1653# a_1419_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u
X36 a_2093_5487# a_591_4917# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X37 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X38 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X39 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X40 vss a_2461_2223# a_393_5042# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 vss a_573_591# a_2461_2223# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X42 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X43 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X44 out1 a_1855_6005# vss vss sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X45 out0 a_1855_6549# vss vss sky130_fd_pr__nfet_01v8 ad=3.51e+11p pd=3.68e+06u as=0p ps=0u w=650000u l=150000u
X46 a_1855_6549# a_2191_6549# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X47 a_591_4917# a_529_6575# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 vss a_529_6575# a_591_4917# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X49 vdd a_843_2741# out4 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X50 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X51 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X52 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X53 vss a_519_4917# a_1179_2741# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X54 vdd a_395_591# a_573_591# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X55 a_841_2223# a_671_2223# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X56 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X57 vdd a_1855_6005# out1 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X58 vdd a_2879_743# a_2879_591# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X59 vss a_697_3311# a_723_3829# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X60 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X61 a_2251_4399# a_1355_1653# a_2191_6549# vdd sky130_fd_pr__pfet_01v8_hvt ad=7.9e+11p pd=7.58e+06u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X62 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X63 vss a_2553_1135# out5 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X64 vss a_519_4917# a_2191_6549# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X65 vdd a_393_5042# a_1635_1653# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X66 vss a_529_6575# a_591_4917# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X67 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X68 vss a_2041_3427# a_2191_6005# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X69 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X70 vdd a_1633_591# out7 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X71 vdd a_529_3311# a_697_3311# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X72 vss a_1633_591# out7 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X73 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X74 a_933_1135# a_763_1135# vss vss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X75 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X76 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X77 out5 a_2553_1135# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X78 out3 a_2879_3855# vss vss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X79 a_1131_1929# a_1355_1653# a_1385_1929# vdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u
X80 vss a_843_2741# out4 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.51e+11p ps=3.68e+06u w=650000u l=150000u
X81 out6 a_2879_591# vss vss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X82 a_2879_743# a_2787_1679# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X83 a_1855_6005# a_2191_6005# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X84 a_1855_6549# a_2191_6549# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X85 out1 a_1855_6005# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X86 out0 a_1855_6549# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X87 a_2431_3311# a_393_5042# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=8.3e+11p pd=7.66e+06u as=0p ps=0u w=1e+06u l=150000u
X88 a_1731_2919# a_573_591# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.5725e+11p pd=2.99e+06u as=0p ps=0u w=420000u l=150000u
X89 vss a_529_3311# a_697_3311# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X90 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X91 vdd a_1131_5495# a_1308_5487# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 a_1225_4399# a_1029_4515# a_1139_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X93 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X94 a_393_5042# a_2461_2223# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X95 out7 a_1633_591# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X96 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X97 vss a_1855_6005# out1 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X98 vss a_1855_6549# out0 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X99 a_2191_6549# a_1355_1653# a_2251_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X100 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X101 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X102 a_573_591# a_395_591# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X103 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X104 a_2879_743# a_2787_1679# vss vss sky130_fd_pr__nfet_01v8 ad=1.352e+11p pd=1.56e+06u as=0p ps=0u w=520000u l=150000u
X105 out5 a_2553_1135# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X106 a_2553_1135# a_841_2223# vss vss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X107 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X108 a_1179_2741# a_1355_1653# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X109 vdd in2 a_395_591# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.65e+11p ps=2.53e+06u w=1e+06u l=150000u
X110 a_1513_2583# a_591_4917# vss vss sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=0p ps=0u w=420000u l=150000u
X111 vss a_529_3311# a_697_3311# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X112 vss a_2553_1135# out5 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X113 vdd a_573_591# a_1636_2455# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.087e+11p ps=1.36e+06u w=420000u l=150000u
X114 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X115 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X116 a_2191_6549# a_1355_1653# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X117 vdd a_749_4943# a_1131_5495# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X118 a_2191_6549# a_393_5042# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X119 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X120 vss a_2093_5487# a_1355_1653# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X121 a_591_4917# a_529_6575# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X122 a_1179_2741# a_1635_1653# a_1385_1929# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X123 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X124 vdd a_841_2223# a_2553_1135# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X125 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X126 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X127 a_749_4943# a_395_4943# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X128 a_2191_6005# a_2041_3427# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X129 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X130 vdd a_697_3311# a_2004_2747# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.087e+11p ps=1.36e+06u w=420000u l=150000u
X131 a_749_4943# a_395_4943# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X132 vdd a_1855_6549# out0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=5.4e+11p ps=5.08e+06u w=1e+06u l=150000u
X133 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X134 a_843_2741# a_1179_2741# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X135 vdd a_723_3829# a_519_4917# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.1e+11p ps=7.62e+06u w=1e+06u l=150000u
X136 vss a_1633_591# out7 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X137 vss a_1855_6005# out1 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X138 vss a_1855_6549# out0 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X139 a_843_2741# a_1179_2741# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X140 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X141 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X142 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X143 vss a_519_4917# a_2191_6005# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X144 a_1633_591# a_1308_5487# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X145 vss a_723_3829# a_519_4917# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5.265e+11p ps=5.52e+06u w=650000u l=150000u
X146 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X147 out3 a_2879_3855# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X148 out4 a_843_2741# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X149 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X150 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X151 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X152 a_1594_2583# a_697_3311# a_1513_2583# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X153 a_1489_1135# a_591_4917# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.087e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X154 out4 a_843_2741# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X155 out1 a_1855_6005# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 vss a_2553_1135# out5 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X157 vss in0 a_529_6575# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X158 vss a_841_2223# a_2553_1135# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X159 a_1355_1653# a_2093_5487# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X160 vss a_1355_1653# a_1179_2741# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X161 a_697_3311# a_529_3311# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X162 vdd a_1355_1653# a_1731_2919# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X163 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X164 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X165 vss a_573_591# a_1748_1495# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X166 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X167 vdd a_763_1367# a_763_1135# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X168 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X169 vss a_1775_4943# out2 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X170 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X171 a_1881_2773# a_573_591# vss vss sky130_fd_pr__nfet_01v8 ad=1.071e+11p pd=1.35e+06u as=0p ps=0u w=420000u l=150000u
X172 vss a_1225_4399# a_1775_4943# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X173 vdd a_2553_1135# out5 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X174 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X175 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X176 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X177 vss a_529_6575# a_591_4917# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X178 a_697_3311# a_529_3311# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X179 a_1179_2741# a_1635_1653# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X180 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X181 vdd a_2553_1135# out5 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X182 out7 a_1633_591# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X183 a_1385_1929# a_1355_1653# a_1131_1929# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X184 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X185 a_393_5042# a_2461_2223# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X186 vdd a_393_5042# a_2431_3311# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X187 vdd a_1225_4399# a_1775_4943# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X188 a_697_3311# a_529_3311# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X189 a_2191_6005# a_2041_3427# a_2151_3311# vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X190 vdd a_573_591# a_1589_1251# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X191 vdd a_519_4917# a_1131_1929# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X192 vss a_2461_2223# a_393_5042# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X193 a_1676_1495# a_1489_1135# a_1589_1251# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.07825e+11p ps=1.36e+06u w=420000u l=150000u
X194 vdd a_723_3829# a_519_4917# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X195 vss a_697_3311# a_2004_2747# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.0785e+11p ps=1.36e+06u w=420000u l=150000u
X196 a_1731_2919# a_2004_2747# a_1962_2773# vss sky130_fd_pr__nfet_01v8 ad=1.07825e+11p pd=1.36e+06u as=8.82e+10p ps=1.26e+06u w=420000u l=150000u
X197 vdd a_1855_6005# out1 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X198 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X199 a_2151_3311# a_519_4917# a_2431_3311# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X200 a_529_3311# in1 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X201 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X202 a_1179_2741# a_519_4917# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X203 vss in1 a_529_3311# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X204 a_2191_6005# a_393_5042# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X205 vdd a_529_6575# a_591_4917# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 a_723_3829# a_697_3311# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X207 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X208 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X209 vss a_573_591# a_1636_2455# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.0785e+11p ps=1.36e+06u w=420000u l=150000u
X210 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X211 out7 a_1633_591# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X212 vss a_1131_5495# a_1308_5487# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X213 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X214 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X215 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X216 a_1731_2919# a_2004_2747# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X217 vss a_843_2741# out4 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X218 a_393_5042# a_2461_2223# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=8.1e+11p pd=7.62e+06u as=0p ps=0u w=1e+06u l=150000u
X219 a_2191_6549# a_519_4917# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X220 out5 a_2553_1135# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X221 a_1029_4515# a_519_4917# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X222 vss a_1775_4943# out2 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X223 vss a_2093_5487# a_1355_1653# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X224 a_591_4917# a_529_6575# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X225 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X226 vss a_2093_5487# a_1355_1653# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X227 vdd a_933_1135# a_2879_3855# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X228 vss a_529_3311# a_697_3311# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X229 out5 a_2553_1135# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X230 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X231 a_723_3829# a_697_3311# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.7e+11p pd=2.54e+06u as=0p ps=0u w=1e+06u l=150000u
X232 a_393_5042# a_2461_2223# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 a_1962_2773# a_1355_1653# a_1881_2773# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X234 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X235 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X236 vdd a_697_3311# a_1363_2455# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.5725e+11p ps=2.99e+06u w=420000u l=150000u
X237 vss a_1308_5487# a_1633_591# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.755e+11p ps=1.84e+06u w=650000u l=150000u
X238 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X239 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X240 a_2553_1135# a_841_2223# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X241 a_393_5042# a_2461_2223# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 a_519_4917# a_723_3829# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X243 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X244 vdd a_393_5042# a_395_4943# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X245 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X246 a_549_4943# a_519_4917# a_477_4943# vss sky130_fd_pr__nfet_01v8 ad=8.82e+10p pd=1.26e+06u as=0p ps=0u w=420000u l=150000u
X247 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X248 out0 a_1855_6549# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X249 vss a_1635_1653# a_1179_2741# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X250 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X251 a_519_4917# a_723_3829# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X252 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X253 vss in2 a_395_591# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X254 vdd a_843_2741# out4 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X255 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X256 vdd a_1775_4943# out2 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X257 vdd a_2879_3855# out3 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X258 a_2041_3427# a_1355_1653# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X259 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X260 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X261 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X262 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X263 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X264 a_2093_5487# a_591_4917# vss vss sky130_fd_pr__nfet_01v8 ad=1.755e+11p pd=1.84e+06u as=0p ps=0u w=650000u l=150000u
X265 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X266 vdd a_393_5042# a_2523_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=8.3e+11p ps=7.66e+06u w=1e+06u l=150000u
X267 out5 a_2553_1135# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X268 a_697_3311# a_529_3311# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X269 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X270 vss a_393_5042# a_2191_6005# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X271 out7 a_1633_591# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X272 vdd a_1633_591# out7 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X273 vdd a_2461_2223# a_393_5042# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X274 vss a_749_4943# a_1131_5495# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X275 vss a_671_2455# a_671_2223# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X276 a_2251_4399# a_519_4917# a_2523_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X277 vss a_1355_1653# a_2191_6549# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X278 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X279 a_1355_1653# a_2093_5487# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X280 vdd a_573_591# a_2461_2223# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.7e+11p ps=2.54e+06u w=1e+06u l=150000u
X281 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X282 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X283 a_1355_1653# a_2093_5487# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X284 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X285 vdd a_529_3311# a_697_3311# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X286 a_1225_4399# a_393_5042# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X287 vdd a_1855_6549# out0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X288 a_1355_1653# a_2093_5487# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X289 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X290 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X291 vss a_1363_2455# a_763_1367# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.69e+11p ps=1.82e+06u w=650000u l=150000u
X292 vss a_393_5042# a_1635_1653# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X293 out4 a_843_2741# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X294 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
X295 out2 a_1775_4943# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X296 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X297 vdd a_529_3311# a_697_3311# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X298 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X299 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X300 out5 a_2553_1135# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X301 a_1131_1929# a_519_4917# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X302 out2 a_1775_4943# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X303 vdd a_1308_5487# a_1633_591# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X304 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X305 a_2431_3311# a_519_4917# a_2151_3311# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X306 a_1225_4399# a_1029_4515# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X307 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X308 a_591_4917# a_529_6575# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X309 vdd in1 a_529_3311# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X310 a_2191_6005# a_519_4917# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X311 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X312 a_519_4917# a_723_3829# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X313 a_2041_3427# a_1355_1653# vss vss sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=0p ps=0u w=420000u l=150000u
X314 a_519_4917# a_723_3829# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X315 out1 a_1855_6005# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X316 a_1363_2455# a_591_4917# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X317 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X318 vdd a_1363_2455# a_763_1367# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.6e+11p ps=2.52e+06u w=1e+06u l=150000u
X319 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X320 a_573_591# a_395_591# vss vss sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=1.38e+06u as=0p ps=0u w=420000u l=150000u
X321 a_933_1135# a_763_1135# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.054e+11p pd=2.1e+06u as=0p ps=0u w=790000u l=150000u
X322 a_1589_1251# a_697_3311# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X323 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X324 a_591_4917# a_529_6575# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X325 vdd a_1633_591# out7 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X326 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X327 a_529_6575# in0 vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X328 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
X329 vss a_591_4917# a_2093_5487# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X330 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X331 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X332 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X333 a_697_3311# a_529_3311# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X334 a_591_4917# a_529_6575# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X335 a_1419_4399# a_393_5042# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X336 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X337 vdd a_2093_5487# a_1355_1653# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X338 vdd a_2553_1135# out5 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X339 vdd a_671_2455# a_671_2223# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X340 a_519_4917# a_723_3829# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X341 a_519_4917# a_723_3829# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X342 vdd a_697_3311# a_723_3829# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X343 vdd a_2461_2223# a_393_5042# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X344 a_1363_2455# a_1636_2455# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X345 a_529_6575# in0 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X346 a_1419_4399# a_1355_1653# a_1139_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X347 vss a_2879_3855# out3 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X348 vdd a_591_4917# a_2093_5487# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X349 out4 a_843_2741# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X350 vdd a_2461_2223# a_393_5042# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X351 vdd a_723_3829# a_519_4917# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X352 vss a_933_1135# a_2879_3855# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X353 a_1945_1135# a_1589_1251# vss vss sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=0p ps=0u w=650000u l=150000u
X354 a_395_4943# a_519_4917# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X355 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X356 vss a_2879_743# a_2879_591# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X357 vss a_393_5042# a_1225_4399# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X358 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X359 a_697_3311# a_529_3311# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X360 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X361 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X362 vss a_2461_2223# a_393_5042# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X363 vss a_2879_591# out6 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X364 vdd a_1945_1135# a_2787_1679# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.054e+11p ps=2.1e+06u w=790000u l=150000u
X365 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X366 vss a_395_591# a_573_591# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X367 vss a_763_1367# a_763_1135# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X368 vss a_1029_4515# a_1225_4399# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X369 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X370 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X371 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X372 a_529_3311# in1 vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X373 a_2151_3311# a_2041_3427# a_2191_6005# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X374 a_2523_4399# a_393_5042# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X375 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X376 vss a_591_4917# a_549_4943# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X377 vss a_1633_591# out7 vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X378 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X379 a_1855_6005# a_2191_6005# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X380 out7 a_1633_591# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X381 out6 a_2879_591# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X382 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
X383 a_1945_1135# a_1589_1251# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=0p ps=0u w=1e+06u l=150000u
X384 a_2523_4399# a_519_4917# a_2251_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X385 a_1308_5487# a_1131_5495# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X386 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
X387 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X388 out2 a_1775_4943# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X389 vdd a_2093_5487# a_1355_1653# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X390 a_1355_1653# a_2093_5487# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X391 vss a_393_5042# a_2191_6549# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X392 a_1225_4399# a_1355_1653# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X393 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X394 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X395 a_1633_591# a_1308_5487# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X396 vss a_1945_1135# a_2787_1679# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.352e+11p ps=1.56e+06u w=520000u l=150000u
X397 vdd a_2093_5487# a_1355_1653# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X398 vss a_723_3829# a_519_4917# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X399 a_2461_2223# a_573_591# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X400 vss a_723_3829# a_519_4917# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X401 vss vdd vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
X402 a_2461_2223# a_573_591# vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X403 vdd vss vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X404 out0 a_1855_6549# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X405 a_1139_4399# a_1029_4515# a_1225_4399# vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

